library verilog;
use verilog.vl_types.all;
entity BCD_seven_seg_A_vlg_vec_tst is
end BCD_seven_seg_A_vlg_vec_tst;
