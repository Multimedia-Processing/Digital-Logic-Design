
`timescale 1ns/1ps

module T;
    reg [7:0] D1 = 8'b01011111;
    reg [7:0] D2 = 8'b01100111;
    wire Eq;


    eq8 UUT (
        .D1(D1),
        .D2(D2),
        .Eq(Eq));
  
    initial
    begin
      #2000 // Final time:  2000 ns
        $stop;
    end

    initial begin
        // -------------  Current Time:  100ns
        #100;
        D1 = 8'b11001000;
        D2 = 8'b10111110;
        // -------------------------------------
        // -------------  Current Time:  200ns
        #100;
        D1 = 8'b10010001;
        D2 = 8'b10010001;
        // -------------------------------------
        // -------------  Current Time:  300ns
        #100;
        D1 = 8'b00011101;
        D2 = 8'b00000101;
        // -------------------------------------
        // -------------  Current Time:  400ns
        #100;
        D1 = 8'b11101010;
        D2 = 8'b11101010;
        // -------------------------------------
        // -------------  Current Time:  500ns
        #100;
        D1 = 8'b01110011;
        D2 = 8'b01011011;
        // -------------------------------------
        // -------------  Current Time:  600ns
        #100;
        D1 = 8'b01110100;
        D2 = 8'b00001111;
        // -------------------------------------
        // -------------  Current Time:  700ns
        #100;
        D1 = 8'b10101000;
        D2 = 8'b10101000;
        // -------------------------------------
        // -------------  Current Time:  800ns
        #100;
        D1 = 8'b00111111;
        D2 = 8'b00011101;
        // -------------------------------------
        // -------------  Current Time:  900ns
        #100;
        D1 = 8'b01100110;
        D2 = 8'b11101110;
        // -------------------------------------
        // -------------  Current Time:  1000ns
        #100;
        D1 = 8'b11001000;
        D2 = 8'b11110010;
        // -------------------------------------
        // -------------  Current Time:  1100ns
        #100;
        D1 = 8'b00011101;
        D2 = 8'b00100101;
        // -------------------------------------
        // -------------  Current Time:  1200ns
        #100;
        D1 = 8'b10000010;
        D2 = 8'b10101100;
        // -------------------------------------
        // -------------  Current Time:  1300ns
        #100;
        D1 = 8'b10000011;
        D2 = 8'b10000011;
        // -------------------------------------
        // -------------  Current Time:  1400ns
        #100;
        D1 = 8'b01011111;
        D2 = 8'b01100111;
        // -------------------------------------
        // -------------  Current Time:  1500ns
        #100;
        D1 = 8'b11001000;
        D2 = 8'b11001000;
        // -------------------------------------
        // -------------  Current Time:  1600ns
        #100;
        D1 = 8'b00100101;
        D2 = 8'b00011001;
        // -------------------------------------
        // -------------  Current Time:  1700ns
        #100;
        D1 = 8'b00111110;
        D2 = 8'b00000101;
        // -------------------------------------
        // -------------  Current Time:  1800ns
        #100;
        D1 = 8'b10101010;
        D2 = 8'b11000010;
        // -------------------------------------
        // -------------  Current Time:  1900ns
        #100;
        D1 = 8'b01100101;
        D2 = 8'b01011111;
        // -------------------------------------
        // -------------  Current Time:  2000ns
        #100;
        D1 = 8'b11110100;
        D2 = 8'b11000100;
    end

endmodule

