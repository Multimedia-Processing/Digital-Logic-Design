module xor_gate(a,b,xor_output);

input a,b;
output xor_output;
xor(xor_output,a,b);

endmodule
