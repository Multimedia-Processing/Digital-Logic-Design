module NAND_GATE (c, a, b);

input a, b;
output c;

    nand(c, a, b);

endmodule 