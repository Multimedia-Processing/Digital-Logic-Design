
`timescale 1ns/1ps

module T;
    reg [3:0] A = 4'b0101;
    reg [3:0] B = 4'b1100;
    reg [3:0] C = 4'b1010;
    reg [3:0] D = 4'b0000;
    reg [1:0] S = 2'b00;
    wire [3:0] Y1;
    wire [3:0] Y2;
    wire [3:0] Y3;


    mux UUT (
        .A(A),
        .B(B),
        .C(C),
        .D(D),
        .S(S),
        .Y1(Y1),
        .Y2(Y2),
        .Y3(Y3));

    initial
    begin
      #2000 // Final time:  2000 ns
        $stop;
    end

    initial begin
        // -------------  Current Time:  100ns
        #100;
        A = 4'b1100;
        B = 4'b1010;
        C = 4'b0011;
        D = 4'b1001;
        // -------------------------------------
        // -------------  Current Time:  200ns
        #100;
        A = 4'b1001;
        B = 4'b0011;
        C = 4'b1111;
        D = 4'b0100;
        // -------------------------------------
        // -------------  Current Time:  300ns
        #100;
        A = 4'b0001;
        B = 4'b1110;
        C = 4'b0100;
        D = 4'b1000;
        // -------------------------------------
        // -------------  Current Time:  400ns
        #100;
        A = 4'b1110;
        B = 4'b0110;
        C = 4'b0101;
        D = 4'b1001;
        // -------------------------------------
        // -------------  Current Time:  500ns
        #100;
        A = 4'b0111;
        B = 4'b0111;
        C = 4'b1001;
        D = 4'b0000;
        S = 2'b01;
        // -------------------------------------
        // -------------  Current Time:  600ns
        #100;
        A = 4'b1001;
        B = 4'b1010;
        C = 4'b0000;
        D = 4'b0010;
        // -------------------------------------
        // -------------  Current Time:  700ns
        #100;
        A = 4'b1010;
        B = 4'b0000;
        C = 4'b0101;
        D = 4'b1111;
        // -------------------------------------
        // -------------  Current Time:  800ns
        #100;
        A = 4'b0011;
        B = 4'b0101;
        C = 4'b1101;
        D = 4'b0110;
        // -------------------------------------
        // -------------  Current Time:  900ns
        #100;
        A = 4'b0110;
        B = 4'b1100;
        C = 4'b0110;
        D = 4'b1010;
        // -------------------------------------
        // -------------  Current Time:  1000ns
        #100;
        A = 4'b1100;
        B = 4'b0101;
        C = 4'b1011;
        D = 4'b1011;
        S = 2'b10;
        // -------------------------------------
        // -------------  Current Time:  1100ns
        #100;
        A = 4'b0001;
        B = 4'b1001;
        C = 4'b1010;
        D = 4'b0010;
        // -------------------------------------
        // -------------  Current Time:  1200ns
        #100;
        A = 4'b1000;
        B = 4'b1000;
        C = 4'b0110;
        D = 4'b1101;
        // -------------------------------------
        // -------------  Current Time:  1300ns
        #100;
        A = 4'b0000;
        B = 4'b0111;
        C = 4'b1111;
        D = 4'b0101;
        // -------------------------------------
        // -------------  Current Time:  1400ns
        #100;
        A = 4'b0101;
        B = 4'b1111;
        C = 4'b0110;
        D = 4'b0000;
        // -------------------------------------
        // -------------  Current Time:  1500ns
        #100;
        A = 4'b1100;
        B = 4'b0110;
        C = 4'b0000;
        D = 4'b1001;
        S = 2'b11;
        // -------------------------------------
        // -------------  Current Time:  1600ns
        #100;
        A = 4'b0010;
        B = 4'b0011;
        C = 4'b1001;
        D = 4'b0101;
        // -------------------------------------
        // -------------  Current Time:  1700ns
        #100;
        A = 4'b0011;
        B = 4'b1011;
        C = 4'b0100;
        D = 4'b1100;
        // -------------------------------------
        // -------------  Current Time:  1800ns
        #100;
        A = 4'b1010;
        B = 4'b0100;
        C = 4'b1100;
        D = 4'b1111;
        // -------------------------------------
        // -------------  Current Time:  1900ns
        #100;
        A = 4'b0110;
        B = 4'b1101;
        C = 4'b1101;
        D = 4'b0011;
        // -------------------------------------
        // -------------  Current Time:  2000ns
        #100;
        A = 4'b1111;
        B = 4'b1001;
        C = 4'b0000;
        D = 4'b1010;
    end
 
endmodule

