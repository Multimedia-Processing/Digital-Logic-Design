
`timescale 1ns/1ps

module T;
    reg [2:0] A = 3'b000;
    wire [1:0] Y;
    wire [1:0] Z;


    casezx UUT (
        .A(A),
        .Y(Y),
        .Z(Z));
    
    initial
    begin 
      #1000 // Final time:  1000 ns
        $stop;
    end

    initial begin
        // -------------  Current Time:  100ns
        #100;
        A = 3'b001;
        // -------------------------------------
        // -------------  Current Time:  200ns
        #100;
        A = 3'b010;
        // -------------------------------------
        // -------------  Current Time:  300ns
        #100;
        A = 3'b011;
        // -------------------------------------
        // -------------  Current Time:  400ns
        #100;
        A = 3'b100;
        // -------------------------------------
        // -------------  Current Time:  500ns
        #100;
        A = 3'b101;
        // -------------------------------------
        // -------------  Current Time:  600ns
        #100;
        A = 3'b110;
        // -------------------------------------
        // -------------  Current Time:  700ns
        #100;
        A = 3'b111;
    end
 
endmodule

