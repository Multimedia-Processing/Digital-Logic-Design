module xnor_gate(a,b,xnor_output);

input a,b;
output xnor_output;
xnor(xnor_output,a,b);

endmodule
