module div_8_assign (a, b, s);
input signed [7:0] a, b;
output signed [8:0] s;

assign s = c / d;

endmodule // div_8_assign
