
`timescale 1ns/1ps

module T;
    reg [3:0] D = 4'b0101;
    wire [3:0] Y1;
    wire [3:0] Y2;
    wire [3:0] Z1;
    wire [3:0] Z2;


    shift_c UUT (
        .D(D),
        .Y1(Y1),
        .Y2(Y2),
        .Z1(Z1),
        .Z2(Z2));

        initial
        begin
          #1000 // Final time:  1000 ns
            $stop;
        end

                initial begin
                    // -------------  Current Time:  100ns
                    #100;
                    D = 4'b1100;
                    // -------------------------------------
                    // -------------  Current Time:  200ns
                    #100;
                    D = 4'b1001;
                    // -------------------------------------
                    // -------------  Current Time:  300ns
                    #100;
                    D = 4'b0001;
                    // -------------------------------------
                    // -------------  Current Time:  400ns
                    #100;
                    D = 4'b1110;
                    // -------------------------------------
                    // -------------  Current Time:  500ns
                    #100;
                    D = 4'b0111;
                    // -------------------------------------
                    // -------------  Current Time:  600ns
                    #100;
                    D = 4'b1001;
                    // -------------------------------------
                    // -------------  Current Time:  700ns
                    #100;
                    D = 4'b1010;
                    // -------------------------------------
                    // -------------  Current Time:  800ns
                    #100;
                    D = 4'b0011;
                    // -------------------------------------
                    // -------------  Current Time:  900ns
                    #100;
                    D = 4'b0110;
                    // -------------------------------------
                    // -------------  Current Time:  1000ns
                    #100;
                    D = 4'b1100;
                end

            endmodule

