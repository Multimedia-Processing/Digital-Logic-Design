module and_gate(a,b,and_output);

input a,b;
output and_output;
and(and_output,a,b);

endmodule
