module xor_gate (a, b, c);

  input a, b ;
  output c ;

  xor (c, a, b);

endmodule // xor_gate
