library verilog;
use verilog.vl_types.all;
entity three_line_to_eight_decimal_decoder_vlg_vec_tst is
end three_line_to_eight_decimal_decoder_vlg_vec_tst;
