// Ch07 adder_4_signed.v
// 四位元有號數加法器

module adder_4_signed ();

endmodule // adder_4_signed
