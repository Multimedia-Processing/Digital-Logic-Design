module or_gate (A,B,C);
    input A,B;
    output C;
    
    or(C,A,B);
    
endmodule