
`timescale 1ns/1ps

module T;
    reg Clk = 1'b0;
    reg Clr = 1'b1;
    reg [1:3] C = 3'b111;
    wire [4:1] R;
    wire [3:0] N;

    parameter PERIOD = 200;
    parameter real DUTY_CYCLE = 0.5;
    parameter OFFSET = 0;

    initial    // Clock process for Clk
    begin
        #OFFSET;
        forever
        begin
            Clk = 1'b0;
            #(PERIOD-(PERIOD*DUTY_CYCLE)) Clk = 1'b1;
            #(PERIOD*DUTY_CYCLE);
        end
    end

    kb1 UUT (
        .Clk(Clk),
        .Clr(Clr),
        .C(C),
        .R(R),
        .N(N));

    initial
    begin
      #4200 // Final time:  4200 ns
        $stop;
    end

    initial begin
        // -------------  Current Time:  115ns
        #115;
        CHECK_N(4'b1111);
        CHECK_R(4'b1110);
        // -------------------------------------
        // -------------  Current Time:  285ns
        #170;
        Clr = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  315ns
        #30;
        CHECK_R(4'b1101);
        // -------------------------------------
        // -------------  Current Time:  515ns
        #200;
        CHECK_R(4'b1011);
        // -------------------------------------
        // -------------  Current Time:  715ns
        #200;
        CHECK_R(4'b0111);
        // -------------------------------------
        // -------------  Current Time:  885ns
        #170;
        C = 3'b011;
        // -------------------------------------
        // -------------  Current Time:  915ns
        #30;
        CHECK_R(4'b1110);
        // -------------------------------------
        // -------------  Current Time:  1115ns
        #200;
        CHECK_R(4'b1101);
        // -------------------------------------
        // -------------  Current Time:  1315ns
        #200;
        CHECK_R(4'b1011);
        // -------------------------------------
        // -------------  Current Time:  1515ns
        #200;
        CHECK_R(4'b0111);
        // -------------------------------------
        // -------------  Current Time:  1685ns
        #170;
        C = 3'b101;
        // -------------------------------------
        // -------------  Current Time:  1715ns
        #30;
        CHECK_R(4'b1110);
        // -------------------------------------
        // -------------  Current Time:  1915ns
        #200;
        CHECK_R(4'b1101);
        // -------------------------------------
        // -------------  Current Time:  2115ns
        #200;
        CHECK_R(4'b1011);
        // -------------------------------------
        // -------------  Current Time:  2315ns
        #200;
        CHECK_R(4'b0111);
        // -------------------------------------
        // -------------  Current Time:  2485ns
        #170;
        C = 3'b110;
        // -------------------------------------
        // -------------  Current Time:  2515ns
        #30;
        CHECK_R(4'b1110);
        // -------------------------------------
        // -------------  Current Time:  2715ns
        #200;
        CHECK_R(4'b1101);
        // -------------------------------------
        // -------------  Current Time:  2915ns
        #200;
        CHECK_R(4'b1011);
        // -------------------------------------
        // -------------  Current Time:  3115ns
        #200;
        CHECK_R(4'b0111);
        // -------------------------------------
        // -------------  Current Time:  3285ns
        #170;
        C = 3'b111;
        // -------------------------------------
        // -------------  Current Time:  3315ns
        #30;
        CHECK_R(4'b1110);
        // -------------------------------------
        // -------------  Current Time:  3515ns
        #200;
        CHECK_R(4'b1101);
        // -------------------------------------
        // -------------  Current Time:  3715ns
        #200;
        CHECK_R(4'b1011);
        // -------------------------------------
        // -------------  Current Time:  3915ns
        #200;
        CHECK_R(4'b0111);
        // -------------------------------------
    end

endmodule

