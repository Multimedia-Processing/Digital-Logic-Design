module xor_gate (a, b, c);
  // 輸入輸出宣告
  input a, b;
  output c;

  // 資料類型宣告
  xor(c, a, b);
    
  // 描述模組內部電路敘述
endmodule // xor_gate