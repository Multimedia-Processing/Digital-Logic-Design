module or_gate(a,b,or_output);

input a,b;
output or_output;
or(or_output,a,b);

endmodule
