// Ch10 kb1.v
// ��L���y��J

module kb1 (Clk, Clr, C, R, N);
input  Clk, Clr;	// �@�줸��J
input  [1:3]  C;	// �T�줸��J
output [4:1]  R;	// �|�줸��X
output [3:0]  N;	// �|�줸��X
reg    [4:1]  R;	// �ŧi���Ȧs�����
reg    [3:0]  N;	// �ŧi���Ȧs�����

// ���ͦ汽�y�H�� R, �`������
always@ (posedge Clk)
  begin
    if (Clr)
      R = 4'b1110;			// R ��� (�u�঳�@��0)
    else
      R = {R[3:1],R[4]};		// �`������

// ����C���, ���䵲�G�s�J N
    case ({R,C})
      7'b1110011  : N = 4'b0001;  	// 1
      7'b1110101  : N = 4'b0010;  	// 2
      7'b1110110  : N = 4'b0011;  	// 3
      7'b1101011  : N = 4'b0100;  	// 4
      7'b1101101  : N = 4'b0101;  	// 5
      7'b1101110  : N = 4'b0110;  	// 6
      7'b1011011  : N = 4'b0111;  	// 7
      7'b1011101  : N = 4'b1000; 	// 8
      7'b1011110  : N = 4'b1001;  	// 9
      7'b0111011  : N = 4'b1010;  	// *
      7'b0111101  : N = 4'b0000;  	// 0
      7'b0111110  : N = 4'b1011;  	// #
      default     : N = N;        	// �����쪬
    endcase
  end

endmodule
