module XOR_GATE (c, a, b);

input a, b;
output c;

    xor(c, a, b);

endmodule