module xnor_gate (A,B,C);
    input A,B;
    output C;
    
    xnor(C,A,B);
    
endmodule