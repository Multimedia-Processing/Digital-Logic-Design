module not_gate (A,C);
    input A;
    output C;
    
    not(C,A);

    
endmodule