
`timescale 1ns/1ps

module T;
    reg [2:0] Q = 3'b000;
    wire [7:0] D1;
    wire [7:0] D2;


    dec38_for_while UUT (
        .Q(Q),
        .D1(D1),
        .D2(D2));

    initial
    begin
      #800 // Final time:  800 ns
        $stop;
    end

    initial begin
        // -------------  Current Time:  100ns
        #100;
        Q = 3'b001;
        // -------------------------------------
        // -------------  Current Time:  200ns
        #100;
        Q = 3'b010;
        // -------------------------------------
        // -------------  Current Time:  300ns
        #100;
        Q = 3'b011;
        // -------------------------------------
        // -------------  Current Time:  400ns
        #100;
        Q = 3'b100;
        // -------------------------------------
        // -------------  Current Time:  500ns
        #100;
        Q = 3'b101;
        // -------------------------------------
        // -------------  Current Time:  600ns
        #100;
        Q = 3'b110;
        // -------------------------------------
        // -------------  Current Time:  700ns
        #100;
        Q = 3'b111;
    end

endmodule

