module nand_gate (A,B,C);
    input A,B;
    output C;
    
    nand(C,A,B);
    
endmodule