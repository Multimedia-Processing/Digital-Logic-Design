`include "full_adder.v"

module full_adder_4_bit ();



endmodule // full_add_4_bit
