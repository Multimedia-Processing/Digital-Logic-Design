module adder_4bit_if(a, b, ci, s, co);
    input [3:0] a,b;
    input ci;
    output [3:0] s;
    output [1:0] co;
    reg [3:0] s;
    reg [1:0] co; 

    always@(a or b or ci)begin
        //  a=0, b=0~F, c=0~1, truth table check ( OK )
        if(         a == 4'b0000 && b == 4'b0000 && ci == 1'b0 )begin     s = 4'b0000;    co = 2'b00;    end
        else if(    a == 4'b0000 && b == 4'b0000 && ci == 1'b1 )begin     s = 4'b0001;    co = 2'b00;    end
        else if(    a == 4'b0000 && b == 4'b0001 && ci == 1'b0 )begin     s = 4'b0001;    co = 2'b00;    end
        else if(    a == 4'b0000 && b == 4'b0001 && ci == 1'b1 )begin     s = 4'b0010;    co = 2'b00;    end
        else if(    a == 4'b0000 && b == 4'b0010 && ci == 1'b0 )begin     s = 4'b0010;    co = 2'b00;    end
        else if(    a == 4'b0000 && b == 4'b0010 && ci == 1'b1 )begin     s = 4'b0011;    co = 2'b00;    end
        else if(    a == 4'b0000 && b == 4'b0011 && ci == 1'b0 )begin     s = 4'b0011;    co = 2'b00;    end
        else if(    a == 4'b0000 && b == 4'b0011 && ci == 1'b1 )begin     s = 4'b0100;    co = 2'b00;    end
        else if(    a == 4'b0000 && b == 4'b0100 && ci == 1'b0 )begin     s = 4'b0100;    co = 2'b00;    end
        else if(    a == 4'b0000 && b == 4'b0100 && ci == 1'b1 )begin     s = 4'b0101;    co = 2'b00;    end
        else if(    a == 4'b0000 && b == 4'b0101 && ci == 1'b0 )begin     s = 4'b0101;    co = 2'b00;    end
        else if(    a == 4'b0000 && b == 4'b0101 && ci == 1'b1 )begin     s = 4'b0110;    co = 2'b00;    end
        else if(    a == 4'b0000 && b == 4'b0110 && ci == 1'b0 )begin     s = 4'b0110;    co = 2'b00;    end
        else if(    a == 4'b0000 && b == 4'b0110 && ci == 1'b1 )begin     s = 4'b0111;    co = 2'b00;    end
        else if(    a == 4'b0000 && b == 4'b0111 && ci == 1'b0 )begin     s = 4'b0111;    co = 2'b00;    end
        else if(    a == 4'b0000 && b == 4'b0111 && ci == 1'b1 )begin     s = 4'b1000;    co = 2'b00;    end
        else if(    a == 4'b0000 && b == 4'b1000 && ci == 1'b0 )begin     s = 4'b1000;    co = 2'b00;    end
        else if(    a == 4'b0000 && b == 4'b1000 && ci == 1'b1 )begin     s = 4'b1001;    co = 2'b00;    end
        else if(    a == 4'b0000 && b == 4'b1001 && ci == 1'b0 )begin     s = 4'b1001;    co = 2'b00;    end
        else if(    a == 4'b0000 && b == 4'b1001 && ci == 1'b1 )begin     s = 4'b1010;    co = 2'b00;    end
        else if(    a == 4'b0000 && b == 4'b1010 && ci == 1'b0 )begin     s = 4'b1010;    co = 2'b00;    end
        else if(    a == 4'b0000 && b == 4'b1010 && ci == 1'b1 )begin     s = 4'b1011;    co = 2'b00;    end
        else if(    a == 4'b0000 && b == 4'b1011 && ci == 1'b0 )begin     s = 4'b1011;    co = 2'b00;    end
        else if(    a == 4'b0000 && b == 4'b1011 && ci == 1'b1 )begin     s = 4'b1100;    co = 2'b00;    end
        else if(    a == 4'b0000 && b == 4'b1100 && ci == 1'b0 )begin     s = 4'b1100;    co = 2'b00;    end
        else if(    a == 4'b0000 && b == 4'b1100 && ci == 1'b1 )begin     s = 4'b1101;    co = 2'b00;    end
        else if(    a == 4'b0000 && b == 4'b1101 && ci == 1'b0 )begin     s = 4'b1101;    co = 2'b00;    end
        else if(    a == 4'b0000 && b == 4'b1101 && ci == 1'b1 )begin     s = 4'b1110;    co = 2'b00;    end
        else if(    a == 4'b0000 && b == 4'b1110 && ci == 1'b0 )begin     s = 4'b1110;    co = 2'b00;    end
        else if(    a == 4'b0000 && b == 4'b1110 && ci == 1'b1 )begin     s = 4'b0000;    co = 2'b01;    end
        else if(    a == 4'b0000 && b == 4'b1111 && ci == 1'b0 )begin     s = 4'b0000;    co = 2'b01;    end
        else if(    a == 4'b0000 && b == 4'b1111 && ci == 1'b1 )begin     s = 4'b0001;    co = 2'b01;    end
        //  a=1, b=0~F, c=0~1, truth table check ( OK )
        else if(    a == 4'b0001 && b == 4'b0000 && ci == 1'b0 )begin     s = 4'b0001;    co = 2'b00;    end
        else if(    a == 4'b0001 && b == 4'b0000 && ci == 1'b1 )begin     s = 4'b0010;    co = 2'b00;    end
        else if(    a == 4'b0001 && b == 4'b0001 && ci == 1'b0 )begin     s = 4'b0010;    co = 2'b00;    end
        else if(    a == 4'b0001 && b == 4'b0001 && ci == 1'b1 )begin     s = 4'b0011;    co = 2'b00;    end
        else if(    a == 4'b0001 && b == 4'b0010 && ci == 1'b0 )begin     s = 4'b0011;    co = 2'b00;    end
        else if(    a == 4'b0001 && b == 4'b0010 && ci == 1'b1 )begin     s = 4'b0100;    co = 2'b00;    end
        else if(    a == 4'b0001 && b == 4'b0011 && ci == 1'b0 )begin     s = 4'b0100;    co = 2'b00;    end
        else if(    a == 4'b0001 && b == 4'b0011 && ci == 1'b1 )begin     s = 4'b0101;    co = 2'b00;    end
        else if(    a == 4'b0001 && b == 4'b0100 && ci == 1'b0 )begin     s = 4'b0101;    co = 2'b00;    end
        else if(    a == 4'b0001 && b == 4'b0100 && ci == 1'b1 )begin     s = 4'b0110;    co = 2'b00;    end
        else if(    a == 4'b0001 && b == 4'b0101 && ci == 1'b0 )begin     s = 4'b0110;    co = 2'b00;    end
        else if(    a == 4'b0001 && b == 4'b0101 && ci == 1'b1 )begin     s = 4'b0111;    co = 2'b00;    end
        else if(    a == 4'b0001 && b == 4'b0110 && ci == 1'b0 )begin     s = 4'b0111;    co = 2'b00;    end
        else if(    a == 4'b0001 && b == 4'b0110 && ci == 1'b1 )begin     s = 4'b1000;    co = 2'b00;    end
        else if(    a == 4'b0001 && b == 4'b0111 && ci == 1'b0 )begin     s = 4'b1000;    co = 2'b00;    end
        else if(    a == 4'b0001 && b == 4'b0111 && ci == 1'b1 )begin     s = 4'b1001;    co = 2'b00;    end
        else if(    a == 4'b0001 && b == 4'b1000 && ci == 1'b0 )begin     s = 4'b1001;    co = 2'b00;    end
        else if(    a == 4'b0001 && b == 4'b1000 && ci == 1'b1 )begin     s = 4'b1010;    co = 2'b00;    end
        else if(    a == 4'b0001 && b == 4'b1001 && ci == 1'b0 )begin     s = 4'b1010;    co = 2'b00;    end
        else if(    a == 4'b0001 && b == 4'b1001 && ci == 1'b1 )begin     s = 4'b1011;    co = 2'b00;    end
        else if(    a == 4'b0001 && b == 4'b1010 && ci == 1'b0 )begin     s = 4'b1011;    co = 2'b00;    end
        else if(    a == 4'b0001 && b == 4'b1010 && ci == 1'b1 )begin     s = 4'b1100;    co = 2'b00;    end
        else if(    a == 4'b0001 && b == 4'b1011 && ci == 1'b0 )begin     s = 4'b1100;    co = 2'b00;    end
        else if(    a == 4'b0001 && b == 4'b1011 && ci == 1'b1 )begin     s = 4'b1101;    co = 2'b00;    end
        else if(    a == 4'b0001 && b == 4'b1100 && ci == 1'b0 )begin     s = 4'b1101;    co = 2'b00;    end
        else if(    a == 4'b0001 && b == 4'b1100 && ci == 1'b1 )begin     s = 4'b1110;    co = 2'b00;    end
        else if(    a == 4'b0001 && b == 4'b1101 && ci == 1'b0 )begin     s = 4'b1110;    co = 2'b00;    end
        else if(    a == 4'b0001 && b == 4'b1101 && ci == 1'b1 )begin     s = 4'b0000;    co = 2'b01;    end
        else if(    a == 4'b0001 && b == 4'b1110 && ci == 1'b0 )begin     s = 4'b0000;    co = 2'b01;    end
        else if(    a == 4'b0001 && b == 4'b1110 && ci == 1'b1 )begin     s = 4'b0001;    co = 2'b01;    end
        else if(    a == 4'b0001 && b == 4'b1111 && ci == 1'b0 )begin     s = 4'b0001;    co = 2'b01;    end
        else if(    a == 4'b0001 && b == 4'b1111 && ci == 1'b1 )begin     s = 4'b0010;    co = 2'b01;    end
        //  a=2, b=0~F, c=0~1, truth table check ( OK )
        else if(    a == 4'b0010 && b == 4'b0000 && ci == 1'b0 )begin     s = 4'b0010;    co = 2'b00;    end
        else if(    a == 4'b0010 && b == 4'b0000 && ci == 1'b1 )begin     s = 4'b0011;    co = 2'b00;    end
        else if(    a == 4'b0010 && b == 4'b0001 && ci == 1'b0 )begin     s = 4'b0011;    co = 2'b00;    end
        else if(    a == 4'b0010 && b == 4'b0001 && ci == 1'b1 )begin     s = 4'b0100;    co = 2'b00;    end
        else if(    a == 4'b0010 && b == 4'b0010 && ci == 1'b0 )begin     s = 4'b0100;    co = 2'b00;    end
        else if(    a == 4'b0010 && b == 4'b0010 && ci == 1'b1 )begin     s = 4'b0101;    co = 2'b00;    end
        else if(    a == 4'b0010 && b == 4'b0011 && ci == 1'b0 )begin     s = 4'b0101;    co = 2'b00;    end
        else if(    a == 4'b0010 && b == 4'b0011 && ci == 1'b1 )begin     s = 4'b0110;    co = 2'b00;    end
        else if(    a == 4'b0010 && b == 4'b0100 && ci == 1'b0 )begin     s = 4'b0110;    co = 2'b00;    end
        else if(    a == 4'b0010 && b == 4'b0100 && ci == 1'b1 )begin     s = 4'b0111;    co = 2'b00;    end
        else if(    a == 4'b0010 && b == 4'b0101 && ci == 1'b0 )begin     s = 4'b0111;    co = 2'b00;    end
        else if(    a == 4'b0010 && b == 4'b0101 && ci == 1'b1 )begin     s = 4'b1000;    co = 2'b00;    end
        else if(    a == 4'b0010 && b == 4'b0110 && ci == 1'b0 )begin     s = 4'b1000;    co = 2'b00;    end
        else if(    a == 4'b0010 && b == 4'b0110 && ci == 1'b1 )begin     s = 4'b1001;    co = 2'b00;    end
        else if(    a == 4'b0010 && b == 4'b0111 && ci == 1'b0 )begin     s = 4'b1001;    co = 2'b00;    end
        else if(    a == 4'b0010 && b == 4'b0111 && ci == 1'b1 )begin     s = 4'b1010;    co = 2'b00;    end
        else if(    a == 4'b0010 && b == 4'b1000 && ci == 1'b0 )begin     s = 4'b1010;    co = 2'b00;    end
        else if(    a == 4'b0010 && b == 4'b1000 && ci == 1'b1 )begin     s = 4'b1011;    co = 2'b00;    end
        else if(    a == 4'b0010 && b == 4'b1001 && ci == 1'b0 )begin     s = 4'b1011;    co = 2'b00;    end
        else if(    a == 4'b0010 && b == 4'b1001 && ci == 1'b1 )begin     s = 4'b1100;    co = 2'b00;    end
        else if(    a == 4'b0010 && b == 4'b1010 && ci == 1'b0 )begin     s = 4'b1100;    co = 2'b00;    end
        else if(    a == 4'b0010 && b == 4'b1010 && ci == 1'b1 )begin     s = 4'b1101;    co = 2'b00;    end
        else if(    a == 4'b0010 && b == 4'b1011 && ci == 1'b0 )begin     s = 4'b1101;    co = 2'b00;    end
        else if(    a == 4'b0010 && b == 4'b1011 && ci == 1'b1 )begin     s = 4'b1110;    co = 2'b00;    end
        else if(    a == 4'b0010 && b == 4'b1100 && ci == 1'b0 )begin     s = 4'b1110;    co = 2'b00;    end
        else if(    a == 4'b0010 && b == 4'b1100 && ci == 1'b1 )begin     s = 4'b0000;    co = 2'b01;    end
        else if(    a == 4'b0010 && b == 4'b1101 && ci == 1'b0 )begin     s = 4'b0000;    co = 2'b01;    end
        else if(    a == 4'b0010 && b == 4'b1101 && ci == 1'b1 )begin     s = 4'b0001;    co = 2'b01;    end
        else if(    a == 4'b0010 && b == 4'b1110 && ci == 1'b0 )begin     s = 4'b0001;    co = 2'b01;    end
        else if(    a == 4'b0010 && b == 4'b1110 && ci == 1'b1 )begin     s = 4'b0010;    co = 2'b01;    end
        else if(    a == 4'b0010 && b == 4'b1111 && ci == 1'b0 )begin     s = 4'b0010;    co = 2'b01;    end
        else if(    a == 4'b0010 && b == 4'b1111 && ci == 1'b1 )begin     s = 4'b0011;    co = 2'b01;    end
        //  a=3, b=0~F, c=0~1, truth table check ( OK )
        else if(    a == 4'b0011 && b == 4'b0000 && ci == 1'b0 )begin     s = 4'b0011;    co = 2'b00;    end
        else if(    a == 4'b0011 && b == 4'b0000 && ci == 1'b1 )begin     s = 4'b0100;    co = 2'b00;    end
        else if(    a == 4'b0011 && b == 4'b0001 && ci == 1'b0 )begin     s = 4'b0100;    co = 2'b00;    end
        else if(    a == 4'b0011 && b == 4'b0001 && ci == 1'b1 )begin     s = 4'b0101;    co = 2'b00;    end
        else if(    a == 4'b0011 && b == 4'b0010 && ci == 1'b0 )begin     s = 4'b0101;    co = 2'b00;    end
        else if(    a == 4'b0011 && b == 4'b0010 && ci == 1'b1 )begin     s = 4'b0110;    co = 2'b00;    end
        else if(    a == 4'b0011 && b == 4'b0011 && ci == 1'b0 )begin     s = 4'b0110;    co = 2'b00;    end
        else if(    a == 4'b0011 && b == 4'b0011 && ci == 1'b1 )begin     s = 4'b0111;    co = 2'b00;    end
        else if(    a == 4'b0011 && b == 4'b0100 && ci == 1'b0 )begin     s = 4'b0111;    co = 2'b00;    end
        else if(    a == 4'b0011 && b == 4'b0100 && ci == 1'b1 )begin     s = 4'b1000;    co = 2'b00;    end
        else if(    a == 4'b0011 && b == 4'b0101 && ci == 1'b0 )begin     s = 4'b1000;    co = 2'b00;    end
        else if(    a == 4'b0011 && b == 4'b0101 && ci == 1'b1 )begin     s = 4'b1001;    co = 2'b00;    end
        else if(    a == 4'b0011 && b == 4'b0110 && ci == 1'b0 )begin     s = 4'b1001;    co = 2'b00;    end
        else if(    a == 4'b0011 && b == 4'b0110 && ci == 1'b1 )begin     s = 4'b1010;    co = 2'b00;    end
        else if(    a == 4'b0011 && b == 4'b0111 && ci == 1'b0 )begin     s = 4'b1010;    co = 2'b00;    end
        else if(    a == 4'b0011 && b == 4'b0111 && ci == 1'b1 )begin     s = 4'b1011;    co = 2'b00;    end
        else if(    a == 4'b0011 && b == 4'b1000 && ci == 1'b0 )begin     s = 4'b1011;    co = 2'b00;    end
        else if(    a == 4'b0011 && b == 4'b1000 && ci == 1'b1 )begin     s = 4'b1100;    co = 2'b00;    end
        else if(    a == 4'b0011 && b == 4'b1001 && ci == 1'b0 )begin     s = 4'b1100;    co = 2'b00;    end
        else if(    a == 4'b0011 && b == 4'b1001 && ci == 1'b1 )begin     s = 4'b1101;    co = 2'b00;    end
        else if(    a == 4'b0011 && b == 4'b1010 && ci == 1'b0 )begin     s = 4'b1101;    co = 2'b00;    end
        else if(    a == 4'b0011 && b == 4'b1010 && ci == 1'b1 )begin     s = 4'b1110;    co = 2'b00;    end
        else if(    a == 4'b0011 && b == 4'b1011 && ci == 1'b0 )begin     s = 4'b1110;    co = 2'b00;    end
        else if(    a == 4'b0011 && b == 4'b1011 && ci == 1'b1 )begin     s = 4'b0000;    co = 2'b01;    end
        else if(    a == 4'b0011 && b == 4'b1100 && ci == 1'b0 )begin     s = 4'b0000;    co = 2'b01;    end
        else if(    a == 4'b0011 && b == 4'b1100 && ci == 1'b1 )begin     s = 4'b0001;    co = 2'b01;    end
        else if(    a == 4'b0011 && b == 4'b1101 && ci == 1'b0 )begin     s = 4'b0001;    co = 2'b01;    end
        else if(    a == 4'b0011 && b == 4'b1101 && ci == 1'b1 )begin     s = 4'b0010;    co = 2'b01;    end
        else if(    a == 4'b0011 && b == 4'b1110 && ci == 1'b0 )begin     s = 4'b0010;    co = 2'b01;    end
        else if(    a == 4'b0011 && b == 4'b1110 && ci == 1'b1 )begin     s = 4'b0011;    co = 2'b01;    end
        else if(    a == 4'b0011 && b == 4'b1111 && ci == 1'b0 )begin     s = 4'b0011;    co = 2'b01;    end
        else if(    a == 4'b0011 && b == 4'b1111 && ci == 1'b1 )begin     s = 4'b0100;    co = 2'b01;    end
        //  a=4, b=0~F, c=0~1, truth table check ( OK )
        else if(    a == 4'b0100 && b == 4'b0000 && ci == 1'b0 )begin     s = 4'b0100;    co = 2'b00;    end
        else if(    a == 4'b0100 && b == 4'b0000 && ci == 1'b1 )begin     s = 4'b0101;    co = 2'b00;    end
        else if(    a == 4'b0100 && b == 4'b0001 && ci == 1'b0 )begin     s = 4'b0101;    co = 2'b00;    end
        else if(    a == 4'b0100 && b == 4'b0001 && ci == 1'b1 )begin     s = 4'b0110;    co = 2'b00;    end
        else if(    a == 4'b0100 && b == 4'b0010 && ci == 1'b0 )begin     s = 4'b0110;    co = 2'b00;    end
        else if(    a == 4'b0100 && b == 4'b0010 && ci == 1'b1 )begin     s = 4'b0111;    co = 2'b00;    end
        else if(    a == 4'b0100 && b == 4'b0011 && ci == 1'b0 )begin     s = 4'b0111;    co = 2'b00;    end
        else if(    a == 4'b0100 && b == 4'b0011 && ci == 1'b1 )begin     s = 4'b1000;    co = 2'b00;    end
        else if(    a == 4'b0100 && b == 4'b0100 && ci == 1'b0 )begin     s = 4'b1000;    co = 2'b00;    end
        else if(    a == 4'b0100 && b == 4'b0100 && ci == 1'b1 )begin     s = 4'b1001;    co = 2'b00;    end
        else if(    a == 4'b0100 && b == 4'b0101 && ci == 1'b0 )begin     s = 4'b1001;    co = 2'b00;    end
        else if(    a == 4'b0100 && b == 4'b0101 && ci == 1'b1 )begin     s = 4'b1010;    co = 2'b00;    end
        else if(    a == 4'b0100 && b == 4'b0110 && ci == 1'b0 )begin     s = 4'b1010;    co = 2'b00;    end
        else if(    a == 4'b0100 && b == 4'b0110 && ci == 1'b1 )begin     s = 4'b1011;    co = 2'b00;    end
        else if(    a == 4'b0100 && b == 4'b0111 && ci == 1'b0 )begin     s = 4'b1011;    co = 2'b00;    end
        else if(    a == 4'b0100 && b == 4'b0111 && ci == 1'b1 )begin     s = 4'b1100;    co = 2'b00;    end
        else if(    a == 4'b0100 && b == 4'b1000 && ci == 1'b0 )begin     s = 4'b1100;    co = 2'b00;    end
        else if(    a == 4'b0100 && b == 4'b1000 && ci == 1'b1 )begin     s = 4'b1101;    co = 2'b00;    end
        else if(    a == 4'b0100 && b == 4'b1001 && ci == 1'b0 )begin     s = 4'b1101;    co = 2'b00;    end
        else if(    a == 4'b0100 && b == 4'b1001 && ci == 1'b1 )begin     s = 4'b1110;    co = 2'b00;    end
        else if(    a == 4'b0100 && b == 4'b1010 && ci == 1'b0 )begin     s = 4'b1110;    co = 2'b00;    end
        else if(    a == 4'b0100 && b == 4'b1010 && ci == 1'b1 )begin     s = 4'b0000;    co = 2'b01;    end
        else if(    a == 4'b0100 && b == 4'b1011 && ci == 1'b0 )begin     s = 4'b0000;    co = 2'b01;    end
        else if(    a == 4'b0100 && b == 4'b1011 && ci == 1'b1 )begin     s = 4'b0001;    co = 2'b01;    end
        else if(    a == 4'b0100 && b == 4'b1100 && ci == 1'b0 )begin     s = 4'b0001;    co = 2'b01;    end
        else if(    a == 4'b0100 && b == 4'b1100 && ci == 1'b1 )begin     s = 4'b0010;    co = 2'b01;    end
        else if(    a == 4'b0100 && b == 4'b1101 && ci == 1'b0 )begin     s = 4'b0010;    co = 2'b01;    end
        else if(    a == 4'b0100 && b == 4'b1101 && ci == 1'b1 )begin     s = 4'b0011;    co = 2'b01;    end
        else if(    a == 4'b0100 && b == 4'b1110 && ci == 1'b0 )begin     s = 4'b0011;    co = 2'b01;    end
        else if(    a == 4'b0100 && b == 4'b1110 && ci == 1'b1 )begin     s = 4'b0100;    co = 2'b01;    end
        else if(    a == 4'b0100 && b == 4'b1111 && ci == 1'b0 )begin     s = 4'b0100;    co = 2'b01;    end
        else if(    a == 4'b0100 && b == 4'b1111 && ci == 1'b1 )begin     s = 4'b0101;    co = 2'b01;    end
        //  a=5, b=0~F, c=0~1, truth table check ( OK )
        else if(    a == 4'b0101 && b == 4'b0000 && ci == 1'b0 )begin     s = 4'b0101;    co = 2'b00;    end
        else if(    a == 4'b0101 && b == 4'b0000 && ci == 1'b1 )begin     s = 4'b0110;    co = 2'b00;    end
        else if(    a == 4'b0101 && b == 4'b0001 && ci == 1'b0 )begin     s = 4'b0110;    co = 2'b00;    end
        else if(    a == 4'b0101 && b == 4'b0001 && ci == 1'b1 )begin     s = 4'b0111;    co = 2'b00;    end
        else if(    a == 4'b0101 && b == 4'b0010 && ci == 1'b0 )begin     s = 4'b0111;    co = 2'b00;    end
        else if(    a == 4'b0101 && b == 4'b0010 && ci == 1'b1 )begin     s = 4'b1000;    co = 2'b00;    end
        else if(    a == 4'b0101 && b == 4'b0011 && ci == 1'b0 )begin     s = 4'b1000;    co = 2'b00;    end
        else if(    a == 4'b0101 && b == 4'b0011 && ci == 1'b1 )begin     s = 4'b1001;    co = 2'b00;    end
        else if(    a == 4'b0101 && b == 4'b0100 && ci == 1'b0 )begin     s = 4'b1001;    co = 2'b00;    end
        else if(    a == 4'b0101 && b == 4'b0100 && ci == 1'b1 )begin     s = 4'b1010;    co = 2'b00;    end
        else if(    a == 4'b0101 && b == 4'b0101 && ci == 1'b0 )begin     s = 4'b1010;    co = 2'b00;    end
        else if(    a == 4'b0101 && b == 4'b0101 && ci == 1'b1 )begin     s = 4'b1011;    co = 2'b00;    end
        else if(    a == 4'b0101 && b == 4'b0110 && ci == 1'b0 )begin     s = 4'b1011;    co = 2'b00;    end
        else if(    a == 4'b0101 && b == 4'b0110 && ci == 1'b1 )begin     s = 4'b1100;    co = 2'b00;    end
        else if(    a == 4'b0101 && b == 4'b0111 && ci == 1'b0 )begin     s = 4'b1100;    co = 2'b00;    end
        else if(    a == 4'b0101 && b == 4'b0111 && ci == 1'b1 )begin     s = 4'b1101;    co = 2'b00;    end
        else if(    a == 4'b0101 && b == 4'b1000 && ci == 1'b0 )begin     s = 4'b1101;    co = 2'b00;    end
        else if(    a == 4'b0101 && b == 4'b1000 && ci == 1'b1 )begin     s = 4'b1110;    co = 2'b00;    end
        else if(    a == 4'b0101 && b == 4'b1001 && ci == 1'b0 )begin     s = 4'b1110;    co = 2'b00;    end
        else if(    a == 4'b0101 && b == 4'b1001 && ci == 1'b1 )begin     s = 4'b0000;    co = 2'b01;    end
        else if(    a == 4'b0101 && b == 4'b1010 && ci == 1'b0 )begin     s = 4'b0000;    co = 2'b01;    end
        else if(    a == 4'b0101 && b == 4'b1010 && ci == 1'b1 )begin     s = 4'b0001;    co = 2'b01;    end
        else if(    a == 4'b0101 && b == 4'b1011 && ci == 1'b0 )begin     s = 4'b0001;    co = 2'b01;    end
        else if(    a == 4'b0101 && b == 4'b1011 && ci == 1'b1 )begin     s = 4'b0010;    co = 2'b01;    end
        else if(    a == 4'b0101 && b == 4'b1100 && ci == 1'b0 )begin     s = 4'b0010;    co = 2'b01;    end
        else if(    a == 4'b0101 && b == 4'b1100 && ci == 1'b1 )begin     s = 4'b0011;    co = 2'b01;    end
        else if(    a == 4'b0101 && b == 4'b1101 && ci == 1'b0 )begin     s = 4'b0011;    co = 2'b01;    end
        else if(    a == 4'b0101 && b == 4'b1101 && ci == 1'b1 )begin     s = 4'b0100;    co = 2'b01;    end
        else if(    a == 4'b0101 && b == 4'b1110 && ci == 1'b0 )begin     s = 4'b0100;    co = 2'b01;    end
        else if(    a == 4'b0101 && b == 4'b1110 && ci == 1'b1 )begin     s = 4'b0101;    co = 2'b01;    end
        else if(    a == 4'b0101 && b == 4'b1111 && ci == 1'b0 )begin     s = 4'b0101;    co = 2'b01;    end
        else if(    a == 4'b0101 && b == 4'b1111 && ci == 1'b1 )begin     s = 4'b0110;    co = 2'b01;    end
        //  a=6, b=0~F, c=0~1, truth table check ( OK )
        else if(    a == 4'b0110 && b == 4'b0000 && ci == 1'b0 )begin     s = 4'b0110;    co = 2'b00;    end
        else if(    a == 4'b0110 && b == 4'b0000 && ci == 1'b1 )begin     s = 4'b0111;    co = 2'b00;    end
        else if(    a == 4'b0110 && b == 4'b0001 && ci == 1'b0 )begin     s = 4'b0111;    co = 2'b00;    end
        else if(    a == 4'b0110 && b == 4'b0001 && ci == 1'b1 )begin     s = 4'b1000;    co = 2'b00;    end
        else if(    a == 4'b0110 && b == 4'b0010 && ci == 1'b0 )begin     s = 4'b1000;    co = 2'b00;    end
        else if(    a == 4'b0110 && b == 4'b0010 && ci == 1'b1 )begin     s = 4'b1001;    co = 2'b00;    end
        else if(    a == 4'b0110 && b == 4'b0011 && ci == 1'b0 )begin     s = 4'b1001;    co = 2'b00;    end
        else if(    a == 4'b0110 && b == 4'b0011 && ci == 1'b1 )begin     s = 4'b1010;    co = 2'b00;    end
        else if(    a == 4'b0110 && b == 4'b0100 && ci == 1'b0 )begin     s = 4'b1010;    co = 2'b00;    end
        else if(    a == 4'b0110 && b == 4'b0100 && ci == 1'b1 )begin     s = 4'b1011;    co = 2'b00;    end
        else if(    a == 4'b0110 && b == 4'b0101 && ci == 1'b0 )begin     s = 4'b1011;    co = 2'b00;    end
        else if(    a == 4'b0110 && b == 4'b0101 && ci == 1'b1 )begin     s = 4'b1100;    co = 2'b00;    end
        else if(    a == 4'b0110 && b == 4'b0110 && ci == 1'b0 )begin     s = 4'b1100;    co = 2'b00;    end
        else if(    a == 4'b0110 && b == 4'b0110 && ci == 1'b1 )begin     s = 4'b1101;    co = 2'b00;    end
        else if(    a == 4'b0110 && b == 4'b0111 && ci == 1'b0 )begin     s = 4'b1101;    co = 2'b00;    end
        else if(    a == 4'b0110 && b == 4'b0111 && ci == 1'b1 )begin     s = 4'b1110;    co = 2'b00;    end
        else if(    a == 4'b0110 && b == 4'b1000 && ci == 1'b0 )begin     s = 4'b1110;    co = 2'b00;    end
        else if(    a == 4'b0110 && b == 4'b1000 && ci == 1'b1 )begin     s = 4'b0000;    co = 2'b01;    end
        else if(    a == 4'b0110 && b == 4'b1001 && ci == 1'b0 )begin     s = 4'b0000;    co = 2'b01;    end
        else if(    a == 4'b0110 && b == 4'b1001 && ci == 1'b1 )begin     s = 4'b0001;    co = 2'b01;    end
        else if(    a == 4'b0110 && b == 4'b1010 && ci == 1'b0 )begin     s = 4'b0001;    co = 2'b01;    end
        else if(    a == 4'b0110 && b == 4'b1010 && ci == 1'b1 )begin     s = 4'b0010;    co = 2'b01;    end
        else if(    a == 4'b0110 && b == 4'b1011 && ci == 1'b0 )begin     s = 4'b0010;    co = 2'b01;    end
        else if(    a == 4'b0110 && b == 4'b1011 && ci == 1'b1 )begin     s = 4'b0011;    co = 2'b01;    end
        else if(    a == 4'b0110 && b == 4'b1100 && ci == 1'b0 )begin     s = 4'b0011;    co = 2'b01;    end
        else if(    a == 4'b0110 && b == 4'b1100 && ci == 1'b1 )begin     s = 4'b0100;    co = 2'b01;    end
        else if(    a == 4'b0110 && b == 4'b1101 && ci == 1'b0 )begin     s = 4'b0100;    co = 2'b01;    end
        else if(    a == 4'b0110 && b == 4'b1101 && ci == 1'b1 )begin     s = 4'b0101;    co = 2'b01;    end
        else if(    a == 4'b0110 && b == 4'b1110 && ci == 1'b0 )begin     s = 4'b0101;    co = 2'b01;    end
        else if(    a == 4'b0110 && b == 4'b1110 && ci == 1'b1 )begin     s = 4'b0110;    co = 2'b01;    end
        else if(    a == 4'b0110 && b == 4'b1111 && ci == 1'b0 )begin     s = 4'b0110;    co = 2'b01;    end
        else if(    a == 4'b0110 && b == 4'b1111 && ci == 1'b1 )begin     s = 4'b0111;    co = 2'b01;    end
        //  a=7, b=0~F, c=0~1, truth table check ( OK )
        else if(    a == 4'b0111 && b == 4'b0000 && ci == 1'b0 )begin     s = 4'b0111;    co = 2'b00;    end
        else if(    a == 4'b0111 && b == 4'b0000 && ci == 1'b1 )begin     s = 4'b1000;    co = 2'b00;    end
        else if(    a == 4'b0111 && b == 4'b0001 && ci == 1'b0 )begin     s = 4'b1000;    co = 2'b00;    end
        else if(    a == 4'b0111 && b == 4'b0001 && ci == 1'b1 )begin     s = 4'b1001;    co = 2'b00;    end
        else if(    a == 4'b0111 && b == 4'b0010 && ci == 1'b0 )begin     s = 4'b1001;    co = 2'b00;    end
        else if(    a == 4'b0111 && b == 4'b0010 && ci == 1'b1 )begin     s = 4'b1010;    co = 2'b00;    end
        else if(    a == 4'b0111 && b == 4'b0011 && ci == 1'b0 )begin     s = 4'b1010;    co = 2'b00;    end
        else if(    a == 4'b0111 && b == 4'b0011 && ci == 1'b1 )begin     s = 4'b1011;    co = 2'b00;    end
        else if(    a == 4'b0111 && b == 4'b0100 && ci == 1'b0 )begin     s = 4'b1011;    co = 2'b00;    end
        else if(    a == 4'b0111 && b == 4'b0100 && ci == 1'b1 )begin     s = 4'b1100;    co = 2'b00;    end
        else if(    a == 4'b0111 && b == 4'b0101 && ci == 1'b0 )begin     s = 4'b1100;    co = 2'b00;    end
        else if(    a == 4'b0111 && b == 4'b0101 && ci == 1'b1 )begin     s = 4'b1101;    co = 2'b00;    end
        else if(    a == 4'b0111 && b == 4'b0110 && ci == 1'b0 )begin     s = 4'b1101;    co = 2'b00;    end
        else if(    a == 4'b0111 && b == 4'b0110 && ci == 1'b1 )begin     s = 4'b1110;    co = 2'b00;    end
        else if(    a == 4'b0111 && b == 4'b0111 && ci == 1'b0 )begin     s = 4'b1110;    co = 2'b00;    end
        else if(    a == 4'b0111 && b == 4'b0111 && ci == 1'b1 )begin     s = 4'b0000;    co = 2'b01;    end
        else if(    a == 4'b0111 && b == 4'b1000 && ci == 1'b0 )begin     s = 4'b0000;    co = 2'b01;    end
        else if(    a == 4'b0111 && b == 4'b1000 && ci == 1'b1 )begin     s = 4'b0001;    co = 2'b01;    end
        else if(    a == 4'b0111 && b == 4'b1001 && ci == 1'b0 )begin     s = 4'b0001;    co = 2'b01;    end
        else if(    a == 4'b0111 && b == 4'b1001 && ci == 1'b1 )begin     s = 4'b0010;    co = 2'b01;    end
        else if(    a == 4'b0111 && b == 4'b1010 && ci == 1'b0 )begin     s = 4'b0010;    co = 2'b01;    end
        else if(    a == 4'b0111 && b == 4'b1010 && ci == 1'b1 )begin     s = 4'b0011;    co = 2'b01;    end
        else if(    a == 4'b0111 && b == 4'b1011 && ci == 1'b0 )begin     s = 4'b0011;    co = 2'b01;    end
        else if(    a == 4'b0111 && b == 4'b1011 && ci == 1'b1 )begin     s = 4'b0100;    co = 2'b01;    end
        else if(    a == 4'b0111 && b == 4'b1100 && ci == 1'b0 )begin     s = 4'b0100;    co = 2'b01;    end
        else if(    a == 4'b0111 && b == 4'b1100 && ci == 1'b1 )begin     s = 4'b0101;    co = 2'b01;    end
        else if(    a == 4'b0111 && b == 4'b1101 && ci == 1'b0 )begin     s = 4'b0101;    co = 2'b01;    end
        else if(    a == 4'b0111 && b == 4'b1101 && ci == 1'b1 )begin     s = 4'b0110;    co = 2'b01;    end
        else if(    a == 4'b0111 && b == 4'b1110 && ci == 1'b0 )begin     s = 4'b0110;    co = 2'b01;    end
        else if(    a == 4'b0111 && b == 4'b1110 && ci == 1'b1 )begin     s = 4'b0111;    co = 2'b01;    end
        else if(    a == 4'b0111 && b == 4'b1111 && ci == 1'b0 )begin     s = 4'b0111;    co = 2'b01;    end
        else if(    a == 4'b0111 && b == 4'b1111 && ci == 1'b1 )begin     s = 4'b1000;    co = 2'b01;    end
        //  a=8, b=0~F, c=0~1, truth table check ( OK )
        else if(    a == 4'b1000 && b == 4'b0000 && ci == 1'b0 )begin     s = 4'b1000;    co = 2'b00;    end
        else if(    a == 4'b1000 && b == 4'b0000 && ci == 1'b1 )begin     s = 4'b1001;    co = 2'b00;    end
        else if(    a == 4'b1000 && b == 4'b0001 && ci == 1'b0 )begin     s = 4'b1001;    co = 2'b00;    end
        else if(    a == 4'b1000 && b == 4'b0001 && ci == 1'b1 )begin     s = 4'b1010;    co = 2'b00;    end
        else if(    a == 4'b1000 && b == 4'b0010 && ci == 1'b0 )begin     s = 4'b1010;    co = 2'b00;    end
        else if(    a == 4'b1000 && b == 4'b0010 && ci == 1'b1 )begin     s = 4'b1011;    co = 2'b00;    end
        else if(    a == 4'b1000 && b == 4'b0011 && ci == 1'b0 )begin     s = 4'b1011;    co = 2'b00;    end
        else if(    a == 4'b1000 && b == 4'b0011 && ci == 1'b1 )begin     s = 4'b1100;    co = 2'b00;    end
        else if(    a == 4'b1000 && b == 4'b0100 && ci == 1'b0 )begin     s = 4'b1100;    co = 2'b00;    end
        else if(    a == 4'b1000 && b == 4'b0100 && ci == 1'b1 )begin     s = 4'b1101;    co = 2'b00;    end
        else if(    a == 4'b1000 && b == 4'b0101 && ci == 1'b0 )begin     s = 4'b1101;    co = 2'b00;    end
        else if(    a == 4'b1000 && b == 4'b0101 && ci == 1'b1 )begin     s = 4'b1110;    co = 2'b00;    end
        else if(    a == 4'b1000 && b == 4'b0110 && ci == 1'b0 )begin     s = 4'b1110;    co = 2'b00;    end
        else if(    a == 4'b1000 && b == 4'b0110 && ci == 1'b1 )begin     s = 4'b0000;    co = 2'b01;    end
        else if(    a == 4'b1000 && b == 4'b0111 && ci == 1'b0 )begin     s = 4'b0000;    co = 2'b01;    end
        else if(    a == 4'b1000 && b == 4'b0111 && ci == 1'b1 )begin     s = 4'b0001;    co = 2'b01;    end
        else if(    a == 4'b1000 && b == 4'b1000 && ci == 1'b0 )begin     s = 4'b0001;    co = 2'b01;    end
        else if(    a == 4'b1000 && b == 4'b1000 && ci == 1'b1 )begin     s = 4'b0010;    co = 2'b01;    end
        else if(    a == 4'b1000 && b == 4'b1001 && ci == 1'b0 )begin     s = 4'b0010;    co = 2'b01;    end
        else if(    a == 4'b1000 && b == 4'b1001 && ci == 1'b1 )begin     s = 4'b0011;    co = 2'b01;    end
        else if(    a == 4'b1000 && b == 4'b1010 && ci == 1'b0 )begin     s = 4'b0011;    co = 2'b01;    end
        else if(    a == 4'b1000 && b == 4'b1010 && ci == 1'b1 )begin     s = 4'b0100;    co = 2'b01;    end
        else if(    a == 4'b1000 && b == 4'b1011 && ci == 1'b0 )begin     s = 4'b0100;    co = 2'b01;    end
        else if(    a == 4'b1000 && b == 4'b1011 && ci == 1'b1 )begin     s = 4'b0101;    co = 2'b01;    end
        else if(    a == 4'b1000 && b == 4'b1100 && ci == 1'b0 )begin     s = 4'b0101;    co = 2'b01;    end
        else if(    a == 4'b1000 && b == 4'b1100 && ci == 1'b1 )begin     s = 4'b0110;    co = 2'b01;    end
        else if(    a == 4'b1000 && b == 4'b1101 && ci == 1'b0 )begin     s = 4'b0110;    co = 2'b01;    end
        else if(    a == 4'b1000 && b == 4'b1101 && ci == 1'b1 )begin     s = 4'b0111;    co = 2'b01;    end
        else if(    a == 4'b1000 && b == 4'b1110 && ci == 1'b0 )begin     s = 4'b0111;    co = 2'b01;    end
        else if(    a == 4'b1000 && b == 4'b1110 && ci == 1'b1 )begin     s = 4'b1000;    co = 2'b01;    end
        else if(    a == 4'b1000 && b == 4'b1111 && ci == 1'b0 )begin     s = 4'b1000;    co = 2'b01;    end
        else if(    a == 4'b1000 && b == 4'b1111 && ci == 1'b1 )begin     s = 4'b1001;    co = 2'b01;    end
        //  a=9, b=0~F, c=0~1, truth table check ( OK )
        else if(    a == 4'b1001 && b == 4'b0000 && ci == 1'b0 )begin     s = 4'b1001;    co = 2'b00;    end
        else if(    a == 4'b1001 && b == 4'b0000 && ci == 1'b1 )begin     s = 4'b1010;    co = 2'b00;    end
        else if(    a == 4'b1001 && b == 4'b0001 && ci == 1'b0 )begin     s = 4'b1010;    co = 2'b00;    end
        else if(    a == 4'b1001 && b == 4'b0001 && ci == 1'b1 )begin     s = 4'b1011;    co = 2'b00;    end
        else if(    a == 4'b1001 && b == 4'b0010 && ci == 1'b0 )begin     s = 4'b1011;    co = 2'b00;    end
        else if(    a == 4'b1001 && b == 4'b0010 && ci == 1'b1 )begin     s = 4'b1100;    co = 2'b00;    end
        else if(    a == 4'b1001 && b == 4'b0011 && ci == 1'b0 )begin     s = 4'b1100;    co = 2'b00;    end
        else if(    a == 4'b1001 && b == 4'b0011 && ci == 1'b1 )begin     s = 4'b1101;    co = 2'b00;    end
        else if(    a == 4'b1001 && b == 4'b0100 && ci == 1'b0 )begin     s = 4'b1101;    co = 2'b00;    end
        else if(    a == 4'b1001 && b == 4'b0100 && ci == 1'b1 )begin     s = 4'b1110;    co = 2'b00;    end
        else if(    a == 4'b1001 && b == 4'b0101 && ci == 1'b0 )begin     s = 4'b1110;    co = 2'b00;    end
        else if(    a == 4'b1001 && b == 4'b0101 && ci == 1'b1 )begin     s = 4'b0000;    co = 2'b01;    end
        else if(    a == 4'b1001 && b == 4'b0110 && ci == 1'b0 )begin     s = 4'b0000;    co = 2'b01;    end
        else if(    a == 4'b1001 && b == 4'b0110 && ci == 1'b1 )begin     s = 4'b0001;    co = 2'b01;    end
        else if(    a == 4'b1001 && b == 4'b0111 && ci == 1'b0 )begin     s = 4'b0001;    co = 2'b01;    end
        else if(    a == 4'b1001 && b == 4'b0111 && ci == 1'b1 )begin     s = 4'b0010;    co = 2'b01;    end
        else if(    a == 4'b1001 && b == 4'b1000 && ci == 1'b0 )begin     s = 4'b0010;    co = 2'b01;    end
        else if(    a == 4'b1001 && b == 4'b1000 && ci == 1'b1 )begin     s = 4'b0011;    co = 2'b01;    end
        else if(    a == 4'b1001 && b == 4'b1001 && ci == 1'b0 )begin     s = 4'b0011;    co = 2'b01;    end
        else if(    a == 4'b1001 && b == 4'b1001 && ci == 1'b1 )begin     s = 4'b0100;    co = 2'b01;    end
        else if(    a == 4'b1001 && b == 4'b1010 && ci == 1'b0 )begin     s = 4'b0100;    co = 2'b01;    end
        else if(    a == 4'b1001 && b == 4'b1010 && ci == 1'b1 )begin     s = 4'b0101;    co = 2'b01;    end
        else if(    a == 4'b1001 && b == 4'b1011 && ci == 1'b0 )begin     s = 4'b0101;    co = 2'b01;    end
        else if(    a == 4'b1001 && b == 4'b1011 && ci == 1'b1 )begin     s = 4'b0110;    co = 2'b01;    end
        else if(    a == 4'b1001 && b == 4'b1100 && ci == 1'b0 )begin     s = 4'b0110;    co = 2'b01;    end
        else if(    a == 4'b1001 && b == 4'b1100 && ci == 1'b1 )begin     s = 4'b0111;    co = 2'b01;    end
        else if(    a == 4'b1001 && b == 4'b1101 && ci == 1'b0 )begin     s = 4'b0111;    co = 2'b01;    end
        else if(    a == 4'b1001 && b == 4'b1101 && ci == 1'b1 )begin     s = 4'b1000;    co = 2'b01;    end
        else if(    a == 4'b1001 && b == 4'b1110 && ci == 1'b0 )begin     s = 4'b1000;    co = 2'b01;    end
        else if(    a == 4'b1001 && b == 4'b1110 && ci == 1'b1 )begin     s = 4'b1001;    co = 2'b01;    end
        else if(    a == 4'b1001 && b == 4'b1111 && ci == 1'b0 )begin     s = 4'b1001;    co = 2'b01;    end
        else if(    a == 4'b1001 && b == 4'b1111 && ci == 1'b1 )begin     s = 4'b1010;    co = 2'b01;    end
        //  a=A, b=0~F, c=0~1, truth table check ( OK )
        else if(    a == 4'b1010 && b == 4'b0000 && ci == 1'b0 )begin     s = 4'b1010;    co = 2'b00;    end
        else if(    a == 4'b1010 && b == 4'b0000 && ci == 1'b1 )begin     s = 4'b1011;    co = 2'b00;    end
        else if(    a == 4'b1010 && b == 4'b0001 && ci == 1'b0 )begin     s = 4'b1011;    co = 2'b00;    end
        else if(    a == 4'b1010 && b == 4'b0001 && ci == 1'b1 )begin     s = 4'b1100;    co = 2'b00;    end
        else if(    a == 4'b1010 && b == 4'b0010 && ci == 1'b0 )begin     s = 4'b1100;    co = 2'b00;    end
        else if(    a == 4'b1010 && b == 4'b0010 && ci == 1'b1 )begin     s = 4'b1101;    co = 2'b00;    end
        else if(    a == 4'b1010 && b == 4'b0011 && ci == 1'b0 )begin     s = 4'b1101;    co = 2'b00;    end
        else if(    a == 4'b1010 && b == 4'b0011 && ci == 1'b1 )begin     s = 4'b1110;    co = 2'b00;    end
        else if(    a == 4'b1010 && b == 4'b0100 && ci == 1'b0 )begin     s = 4'b1110;    co = 2'b00;    end
        else if(    a == 4'b1010 && b == 4'b0100 && ci == 1'b1 )begin     s = 4'b0000;    co = 2'b01;    end
        else if(    a == 4'b1010 && b == 4'b0101 && ci == 1'b0 )begin     s = 4'b0000;    co = 2'b01;    end
        else if(    a == 4'b1010 && b == 4'b0101 && ci == 1'b1 )begin     s = 4'b0001;    co = 2'b01;    end
        else if(    a == 4'b1010 && b == 4'b0110 && ci == 1'b0 )begin     s = 4'b0001;    co = 2'b01;    end
        else if(    a == 4'b1010 && b == 4'b0110 && ci == 1'b1 )begin     s = 4'b0010;    co = 2'b01;    end
        else if(    a == 4'b1010 && b == 4'b0111 && ci == 1'b0 )begin     s = 4'b0010;    co = 2'b01;    end
        else if(    a == 4'b1010 && b == 4'b0111 && ci == 1'b1 )begin     s = 4'b0011;    co = 2'b01;    end
        else if(    a == 4'b1010 && b == 4'b1000 && ci == 1'b0 )begin     s = 4'b0011;    co = 2'b01;    end
        else if(    a == 4'b1010 && b == 4'b1000 && ci == 1'b1 )begin     s = 4'b0100;    co = 2'b01;    end
        else if(    a == 4'b1010 && b == 4'b1001 && ci == 1'b0 )begin     s = 4'b0100;    co = 2'b01;    end
        else if(    a == 4'b1010 && b == 4'b1001 && ci == 1'b1 )begin     s = 4'b0101;    co = 2'b01;    end
        else if(    a == 4'b1010 && b == 4'b1010 && ci == 1'b0 )begin     s = 4'b0101;    co = 2'b01;    end
        else if(    a == 4'b1010 && b == 4'b1010 && ci == 1'b1 )begin     s = 4'b0110;    co = 2'b01;    end
        else if(    a == 4'b1010 && b == 4'b1011 && ci == 1'b0 )begin     s = 4'b0110;    co = 2'b01;    end
        else if(    a == 4'b1010 && b == 4'b1011 && ci == 1'b1 )begin     s = 4'b0111;    co = 2'b01;    end
        else if(    a == 4'b1010 && b == 4'b1100 && ci == 1'b0 )begin     s = 4'b0111;    co = 2'b01;    end
        else if(    a == 4'b1010 && b == 4'b1100 && ci == 1'b1 )begin     s = 4'b1000;    co = 2'b01;    end
        else if(    a == 4'b1010 && b == 4'b1101 && ci == 1'b0 )begin     s = 4'b1000;    co = 2'b01;    end
        else if(    a == 4'b1010 && b == 4'b1101 && ci == 1'b1 )begin     s = 4'b1001;    co = 2'b01;    end
        else if(    a == 4'b1010 && b == 4'b1110 && ci == 1'b0 )begin     s = 4'b1001;    co = 2'b01;    end
        else if(    a == 4'b1010 && b == 4'b1110 && ci == 1'b1 )begin     s = 4'b1010;    co = 2'b01;    end
        else if(    a == 4'b1010 && b == 4'b1111 && ci == 1'b0 )begin     s = 4'b1010;    co = 2'b01;    end
        else if(    a == 4'b1010 && b == 4'b1111 && ci == 1'b1 )begin     s = 4'b1011;    co = 2'b01;    end
        //  a=B, b=0~F, c=0~1, truth table check ( OK )
        else if(    a == 4'b1011 && b == 4'b0000 && ci == 1'b0 )begin     s = 4'b1011;    co = 2'b00;    end
        else if(    a == 4'b1011 && b == 4'b0000 && ci == 1'b1 )begin     s = 4'b1100;    co = 2'b00;    end
        else if(    a == 4'b1011 && b == 4'b0001 && ci == 1'b0 )begin     s = 4'b1100;    co = 2'b00;    end
        else if(    a == 4'b1011 && b == 4'b0001 && ci == 1'b1 )begin     s = 4'b1101;    co = 2'b00;    end
        else if(    a == 4'b1011 && b == 4'b0010 && ci == 1'b0 )begin     s = 4'b1101;    co = 2'b00;    end
        else if(    a == 4'b1011 && b == 4'b0010 && ci == 1'b1 )begin     s = 4'b1110;    co = 2'b00;    end
        else if(    a == 4'b1011 && b == 4'b0011 && ci == 1'b0 )begin     s = 4'b1110;    co = 2'b00;    end
        else if(    a == 4'b1011 && b == 4'b0011 && ci == 1'b1 )begin     s = 4'b0000;    co = 2'b01;    end
        else if(    a == 4'b1011 && b == 4'b0100 && ci == 1'b0 )begin     s = 4'b0000;    co = 2'b01;    end
        else if(    a == 4'b1011 && b == 4'b0100 && ci == 1'b1 )begin     s = 4'b0001;    co = 2'b01;    end
        else if(    a == 4'b1011 && b == 4'b0101 && ci == 1'b0 )begin     s = 4'b0001;    co = 2'b01;    end
        else if(    a == 4'b1011 && b == 4'b0101 && ci == 1'b1 )begin     s = 4'b0010;    co = 2'b01;    end
        else if(    a == 4'b1011 && b == 4'b0110 && ci == 1'b0 )begin     s = 4'b0010;    co = 2'b01;    end
        else if(    a == 4'b1011 && b == 4'b0110 && ci == 1'b1 )begin     s = 4'b0011;    co = 2'b01;    end
        else if(    a == 4'b1011 && b == 4'b0111 && ci == 1'b0 )begin     s = 4'b0011;    co = 2'b01;    end
        else if(    a == 4'b1011 && b == 4'b0111 && ci == 1'b1 )begin     s = 4'b0100;    co = 2'b01;    end
        else if(    a == 4'b1011 && b == 4'b1000 && ci == 1'b0 )begin     s = 4'b0100;    co = 2'b01;    end
        else if(    a == 4'b1011 && b == 4'b1000 && ci == 1'b1 )begin     s = 4'b0101;    co = 2'b01;    end
        else if(    a == 4'b1011 && b == 4'b1001 && ci == 1'b0 )begin     s = 4'b0101;    co = 2'b01;    end
        else if(    a == 4'b1011 && b == 4'b1001 && ci == 1'b1 )begin     s = 4'b0110;    co = 2'b01;    end
        else if(    a == 4'b1011 && b == 4'b1010 && ci == 1'b0 )begin     s = 4'b0110;    co = 2'b01;    end
        else if(    a == 4'b1011 && b == 4'b1010 && ci == 1'b1 )begin     s = 4'b0111;    co = 2'b01;    end
        else if(    a == 4'b1011 && b == 4'b1011 && ci == 1'b0 )begin     s = 4'b0111;    co = 2'b01;    end
        else if(    a == 4'b1011 && b == 4'b1011 && ci == 1'b1 )begin     s = 4'b1000;    co = 2'b01;    end
        else if(    a == 4'b1011 && b == 4'b1100 && ci == 1'b0 )begin     s = 4'b1000;    co = 2'b01;    end
        else if(    a == 4'b1011 && b == 4'b1100 && ci == 1'b1 )begin     s = 4'b1001;    co = 2'b01;    end
        else if(    a == 4'b1011 && b == 4'b1101 && ci == 1'b0 )begin     s = 4'b1001;    co = 2'b01;    end
        else if(    a == 4'b1011 && b == 4'b1101 && ci == 1'b1 )begin     s = 4'b1010;    co = 2'b01;    end
        else if(    a == 4'b1011 && b == 4'b1110 && ci == 1'b0 )begin     s = 4'b1010;    co = 2'b01;    end
        else if(    a == 4'b1011 && b == 4'b1110 && ci == 1'b1 )begin     s = 4'b1011;    co = 2'b01;    end
        else if(    a == 4'b1011 && b == 4'b1111 && ci == 1'b0 )begin     s = 4'b1011;    co = 2'b01;    end
        else if(    a == 4'b1011 && b == 4'b1111 && ci == 1'b1 )begin     s = 4'b1100;    co = 2'b01;    end
        //  a=C, b=0~F, c=0~1, truth table check ( OK )
        else if(    a == 4'b1100 && b == 4'b0000 && ci == 1'b0 )begin     s = 4'b1100;    co = 2'b00;    end
        else if(    a == 4'b1100 && b == 4'b0000 && ci == 1'b1 )begin     s = 4'b1101;    co = 2'b00;    end
        else if(    a == 4'b1100 && b == 4'b0001 && ci == 1'b0 )begin     s = 4'b1101;    co = 2'b00;    end
        else if(    a == 4'b1100 && b == 4'b0001 && ci == 1'b1 )begin     s = 4'b1110;    co = 2'b00;    end
        else if(    a == 4'b1100 && b == 4'b0010 && ci == 1'b0 )begin     s = 4'b1110;    co = 2'b00;    end
        else if(    a == 4'b1100 && b == 4'b0010 && ci == 1'b1 )begin     s = 4'b0000;    co = 2'b01;    end
        else if(    a == 4'b1100 && b == 4'b0011 && ci == 1'b0 )begin     s = 4'b0000;    co = 2'b01;    end
        else if(    a == 4'b1100 && b == 4'b0011 && ci == 1'b1 )begin     s = 4'b0001;    co = 2'b01;    end
        else if(    a == 4'b1100 && b == 4'b0100 && ci == 1'b0 )begin     s = 4'b0001;    co = 2'b01;    end
        else if(    a == 4'b1100 && b == 4'b0100 && ci == 1'b1 )begin     s = 4'b0010;    co = 2'b01;    end
        else if(    a == 4'b1100 && b == 4'b0101 && ci == 1'b0 )begin     s = 4'b0010;    co = 2'b01;    end
        else if(    a == 4'b1100 && b == 4'b0101 && ci == 1'b1 )begin     s = 4'b0011;    co = 2'b01;    end
        else if(    a == 4'b1100 && b == 4'b0110 && ci == 1'b0 )begin     s = 4'b0011;    co = 2'b01;    end
        else if(    a == 4'b1100 && b == 4'b0110 && ci == 1'b1 )begin     s = 4'b0100;    co = 2'b01;    end
        else if(    a == 4'b1100 && b == 4'b0111 && ci == 1'b0 )begin     s = 4'b0100;    co = 2'b01;    end
        else if(    a == 4'b1100 && b == 4'b0111 && ci == 1'b1 )begin     s = 4'b0101;    co = 2'b01;    end
        else if(    a == 4'b1100 && b == 4'b1000 && ci == 1'b0 )begin     s = 4'b0101;    co = 2'b01;    end
        else if(    a == 4'b1100 && b == 4'b1000 && ci == 1'b1 )begin     s = 4'b0110;    co = 2'b01;    end
        else if(    a == 4'b1100 && b == 4'b1001 && ci == 1'b0 )begin     s = 4'b0110;    co = 2'b01;    end
        else if(    a == 4'b1100 && b == 4'b1001 && ci == 1'b1 )begin     s = 4'b0111;    co = 2'b01;    end
        else if(    a == 4'b1100 && b == 4'b1010 && ci == 1'b0 )begin     s = 4'b0111;    co = 2'b01;    end
        else if(    a == 4'b1100 && b == 4'b1010 && ci == 1'b1 )begin     s = 4'b1000;    co = 2'b01;    end
        else if(    a == 4'b1100 && b == 4'b1011 && ci == 1'b0 )begin     s = 4'b1000;    co = 2'b01;    end
        else if(    a == 4'b1100 && b == 4'b1011 && ci == 1'b1 )begin     s = 4'b1001;    co = 2'b01;    end
        else if(    a == 4'b1100 && b == 4'b1100 && ci == 1'b0 )begin     s = 4'b1001;    co = 2'b01;    end
        else if(    a == 4'b1100 && b == 4'b1100 && ci == 1'b1 )begin     s = 4'b1010;    co = 2'b01;    end
        else if(    a == 4'b1100 && b == 4'b1101 && ci == 1'b0 )begin     s = 4'b1010;    co = 2'b01;    end
        else if(    a == 4'b1100 && b == 4'b1101 && ci == 1'b1 )begin     s = 4'b1011;    co = 2'b01;    end
        else if(    a == 4'b1100 && b == 4'b1110 && ci == 1'b0 )begin     s = 4'b1011;    co = 2'b01;    end
        else if(    a == 4'b1100 && b == 4'b1110 && ci == 1'b1 )begin     s = 4'b1100;    co = 2'b01;    end
        else if(    a == 4'b1100 && b == 4'b1111 && ci == 1'b0 )begin     s = 4'b1100;    co = 2'b01;    end
        else if(    a == 4'b1100 && b == 4'b1111 && ci == 1'b1 )begin     s = 4'b1101;    co = 2'b01;    end
        //  a=D, b=0~F, c=0~1, truth table check ( OK )
        else if(    a == 4'b1101 && b == 4'b0000 && ci == 1'b0 )begin     s = 4'b1101;    co = 2'b00;    end
        else if(    a == 4'b1101 && b == 4'b0000 && ci == 1'b1 )begin     s = 4'b1110;    co = 2'b00;    end
        else if(    a == 4'b1101 && b == 4'b0001 && ci == 1'b0 )begin     s = 4'b1110;    co = 2'b00;    end
        else if(    a == 4'b1101 && b == 4'b0001 && ci == 1'b1 )begin     s = 4'b0000;    co = 2'b01;    end
        else if(    a == 4'b1101 && b == 4'b0010 && ci == 1'b0 )begin     s = 4'b0000;    co = 2'b01;    end
        else if(    a == 4'b1101 && b == 4'b0010 && ci == 1'b1 )begin     s = 4'b0001;    co = 2'b01;    end
        else if(    a == 4'b1101 && b == 4'b0011 && ci == 1'b0 )begin     s = 4'b0001;    co = 2'b01;    end
        else if(    a == 4'b1101 && b == 4'b0011 && ci == 1'b1 )begin     s = 4'b0010;    co = 2'b01;    end
        else if(    a == 4'b1101 && b == 4'b0100 && ci == 1'b0 )begin     s = 4'b0010;    co = 2'b01;    end
        else if(    a == 4'b1101 && b == 4'b0100 && ci == 1'b1 )begin     s = 4'b0011;    co = 2'b01;    end
        else if(    a == 4'b1101 && b == 4'b0101 && ci == 1'b0 )begin     s = 4'b0011;    co = 2'b01;    end
        else if(    a == 4'b1101 && b == 4'b0101 && ci == 1'b1 )begin     s = 4'b0100;    co = 2'b01;    end
        else if(    a == 4'b1101 && b == 4'b0110 && ci == 1'b0 )begin     s = 4'b0100;    co = 2'b01;    end
        else if(    a == 4'b1101 && b == 4'b0110 && ci == 1'b1 )begin     s = 4'b0101;    co = 2'b01;    end
        else if(    a == 4'b1101 && b == 4'b0111 && ci == 1'b0 )begin     s = 4'b0101;    co = 2'b01;    end
        else if(    a == 4'b1101 && b == 4'b0111 && ci == 1'b1 )begin     s = 4'b0110;    co = 2'b01;    end
        else if(    a == 4'b1101 && b == 4'b1000 && ci == 1'b0 )begin     s = 4'b0110;    co = 2'b01;    end
        else if(    a == 4'b1101 && b == 4'b1000 && ci == 1'b1 )begin     s = 4'b0111;    co = 2'b01;    end
        else if(    a == 4'b1101 && b == 4'b1001 && ci == 1'b0 )begin     s = 4'b0111;    co = 2'b01;    end
        else if(    a == 4'b1101 && b == 4'b1001 && ci == 1'b1 )begin     s = 4'b1000;    co = 2'b01;    end
        else if(    a == 4'b1101 && b == 4'b1010 && ci == 1'b0 )begin     s = 4'b1000;    co = 2'b01;    end
        else if(    a == 4'b1101 && b == 4'b1010 && ci == 1'b1 )begin     s = 4'b1001;    co = 2'b01;    end
        else if(    a == 4'b1101 && b == 4'b1011 && ci == 1'b0 )begin     s = 4'b1001;    co = 2'b01;    end
        else if(    a == 4'b1101 && b == 4'b1011 && ci == 1'b1 )begin     s = 4'b1010;    co = 2'b01;    end
        else if(    a == 4'b1101 && b == 4'b1100 && ci == 1'b0 )begin     s = 4'b1010;    co = 2'b01;    end
        else if(    a == 4'b1101 && b == 4'b1100 && ci == 1'b1 )begin     s = 4'b1011;    co = 2'b01;    end
        else if(    a == 4'b1101 && b == 4'b1101 && ci == 1'b0 )begin     s = 4'b1011;    co = 2'b01;    end
        else if(    a == 4'b1101 && b == 4'b1101 && ci == 1'b1 )begin     s = 4'b1100;    co = 2'b01;    end
        else if(    a == 4'b1101 && b == 4'b1110 && ci == 1'b0 )begin     s = 4'b1100;    co = 2'b01;    end
        else if(    a == 4'b1101 && b == 4'b1110 && ci == 1'b1 )begin     s = 4'b1101;    co = 2'b01;    end
        else if(    a == 4'b1101 && b == 4'b1111 && ci == 1'b0 )begin     s = 4'b1101;    co = 2'b01;    end
        else if(    a == 4'b1101 && b == 4'b1111 && ci == 1'b1 )begin     s = 4'b1110;    co = 2'b01;    end
        //  a=E, b=0~F, c=0~1, truth table check ( OK )
        else if(    a == 4'b1110 && b == 4'b0000 && ci == 1'b0 )begin     s = 4'b1110;    co = 2'b00;    end
        else if(    a == 4'b1110 && b == 4'b0000 && ci == 1'b1 )begin     s = 4'b0000;    co = 2'b01;    end
        else if(    a == 4'b1110 && b == 4'b0001 && ci == 1'b0 )begin     s = 4'b0000;    co = 2'b01;    end
        else if(    a == 4'b1110 && b == 4'b0001 && ci == 1'b1 )begin     s = 4'b0001;    co = 2'b01;    end
        else if(    a == 4'b1110 && b == 4'b0010 && ci == 1'b0 )begin     s = 4'b0001;    co = 2'b01;    end
        else if(    a == 4'b1110 && b == 4'b0010 && ci == 1'b1 )begin     s = 4'b0010;    co = 2'b01;    end
        else if(    a == 4'b1110 && b == 4'b0011 && ci == 1'b0 )begin     s = 4'b0010;    co = 2'b01;    end
        else if(    a == 4'b1110 && b == 4'b0011 && ci == 1'b1 )begin     s = 4'b0011;    co = 2'b01;    end
        else if(    a == 4'b1110 && b == 4'b0100 && ci == 1'b0 )begin     s = 4'b0011;    co = 2'b01;    end
        else if(    a == 4'b1110 && b == 4'b0100 && ci == 1'b1 )begin     s = 4'b0100;    co = 2'b01;    end
        else if(    a == 4'b1110 && b == 4'b0101 && ci == 1'b0 )begin     s = 4'b0100;    co = 2'b01;    end
        else if(    a == 4'b1110 && b == 4'b0101 && ci == 1'b1 )begin     s = 4'b0101;    co = 2'b01;    end
        else if(    a == 4'b1110 && b == 4'b0110 && ci == 1'b0 )begin     s = 4'b0101;    co = 2'b01;    end
        else if(    a == 4'b1110 && b == 4'b0110 && ci == 1'b1 )begin     s = 4'b0110;    co = 2'b01;    end
        else if(    a == 4'b1110 && b == 4'b0111 && ci == 1'b0 )begin     s = 4'b0110;    co = 2'b01;    end
        else if(    a == 4'b1110 && b == 4'b0111 && ci == 1'b1 )begin     s = 4'b0111;    co = 2'b01;    end
        else if(    a == 4'b1110 && b == 4'b1000 && ci == 1'b0 )begin     s = 4'b0111;    co = 2'b01;    end
        else if(    a == 4'b1110 && b == 4'b1000 && ci == 1'b1 )begin     s = 4'b1000;    co = 2'b01;    end
        else if(    a == 4'b1110 && b == 4'b1001 && ci == 1'b0 )begin     s = 4'b1000;    co = 2'b01;    end
        else if(    a == 4'b1110 && b == 4'b1001 && ci == 1'b1 )begin     s = 4'b1001;    co = 2'b01;    end
        else if(    a == 4'b1110 && b == 4'b1010 && ci == 1'b0 )begin     s = 4'b1001;    co = 2'b01;    end
        else if(    a == 4'b1110 && b == 4'b1010 && ci == 1'b1 )begin     s = 4'b1010;    co = 2'b01;    end
        else if(    a == 4'b1110 && b == 4'b1011 && ci == 1'b0 )begin     s = 4'b1010;    co = 2'b01;    end
        else if(    a == 4'b1110 && b == 4'b1011 && ci == 1'b1 )begin     s = 4'b1011;    co = 2'b01;    end
        else if(    a == 4'b1110 && b == 4'b1100 && ci == 1'b0 )begin     s = 4'b1011;    co = 2'b01;    end
        else if(    a == 4'b1110 && b == 4'b1100 && ci == 1'b1 )begin     s = 4'b1100;    co = 2'b01;    end
        else if(    a == 4'b1110 && b == 4'b1101 && ci == 1'b0 )begin     s = 4'b1100;    co = 2'b01;    end
        else if(    a == 4'b1110 && b == 4'b1101 && ci == 1'b1 )begin     s = 4'b1101;    co = 2'b01;    end
        else if(    a == 4'b1110 && b == 4'b1110 && ci == 1'b0 )begin     s = 4'b1101;    co = 2'b01;    end
        else if(    a == 4'b1110 && b == 4'b1110 && ci == 1'b1 )begin     s = 4'b1110;    co = 2'b01;    end
        else if(    a == 4'b1110 && b == 4'b1111 && ci == 1'b0 )begin     s = 4'b1110;    co = 2'b01;    end
        else if(    a == 4'b1110 && b == 4'b1111 && ci == 1'b1 )begin     s = 4'b0000;    co = 2'b10;    end
        //  a=F, b=0~F, c=0~1, truth table check ( OK )
        else if(    a == 4'b1111 && b == 4'b0000 && ci == 1'b0 )begin     s = 4'b0000;    co = 2'b01;    end
        else if(    a == 4'b1111 && b == 4'b0000 && ci == 1'b1 )begin     s = 4'b0001;    co = 2'b01;    end
        else if(    a == 4'b1111 && b == 4'b0001 && ci == 1'b0 )begin     s = 4'b0001;    co = 2'b01;    end
        else if(    a == 4'b1111 && b == 4'b0001 && ci == 1'b1 )begin     s = 4'b0010;    co = 2'b01;    end
        else if(    a == 4'b1111 && b == 4'b0010 && ci == 1'b0 )begin     s = 4'b0010;    co = 2'b01;    end
        else if(    a == 4'b1111 && b == 4'b0010 && ci == 1'b1 )begin     s = 4'b0011;    co = 2'b01;    end
        else if(    a == 4'b1111 && b == 4'b0011 && ci == 1'b0 )begin     s = 4'b0011;    co = 2'b01;    end
        else if(    a == 4'b1111 && b == 4'b0011 && ci == 1'b1 )begin     s = 4'b0100;    co = 2'b01;    end
        else if(    a == 4'b1111 && b == 4'b0100 && ci == 1'b0 )begin     s = 4'b0100;    co = 2'b01;    end
        else if(    a == 4'b1111 && b == 4'b0100 && ci == 1'b1 )begin     s = 4'b0101;    co = 2'b01;    end
        else if(    a == 4'b1111 && b == 4'b0101 && ci == 1'b0 )begin     s = 4'b0101;    co = 2'b01;    end
        else if(    a == 4'b1111 && b == 4'b0101 && ci == 1'b1 )begin     s = 4'b0110;    co = 2'b01;    end
        else if(    a == 4'b1111 && b == 4'b0110 && ci == 1'b0 )begin     s = 4'b0110;    co = 2'b01;    end
        else if(    a == 4'b1111 && b == 4'b0110 && ci == 1'b1 )begin     s = 4'b0111;    co = 2'b01;    end
        else if(    a == 4'b1111 && b == 4'b0111 && ci == 1'b0 )begin     s = 4'b0111;    co = 2'b01;    end
        else if(    a == 4'b1111 && b == 4'b0111 && ci == 1'b1 )begin     s = 4'b1000;    co = 2'b01;    end
        else if(    a == 4'b1111 && b == 4'b1000 && ci == 1'b0 )begin     s = 4'b1000;    co = 2'b01;    end
        else if(    a == 4'b1111 && b == 4'b1000 && ci == 1'b1 )begin     s = 4'b1001;    co = 2'b01;    end
        else if(    a == 4'b1111 && b == 4'b1001 && ci == 1'b0 )begin     s = 4'b1001;    co = 2'b01;    end
        else if(    a == 4'b1111 && b == 4'b1001 && ci == 1'b1 )begin     s = 4'b1010;    co = 2'b01;    end
        else if(    a == 4'b1111 && b == 4'b1010 && ci == 1'b0 )begin     s = 4'b1010;    co = 2'b01;    end
        else if(    a == 4'b1111 && b == 4'b1010 && ci == 1'b1 )begin     s = 4'b1011;    co = 2'b01;    end
        else if(    a == 4'b1111 && b == 4'b1011 && ci == 1'b0 )begin     s = 4'b1011;    co = 2'b01;    end
        else if(    a == 4'b1111 && b == 4'b1011 && ci == 1'b1 )begin     s = 4'b1100;    co = 2'b01;    end
        else if(    a == 4'b1111 && b == 4'b1100 && ci == 1'b0 )begin     s = 4'b1100;    co = 2'b01;    end
        else if(    a == 4'b1111 && b == 4'b1100 && ci == 1'b1 )begin     s = 4'b1101;    co = 2'b01;    end
        else if(    a == 4'b1111 && b == 4'b1101 && ci == 1'b0 )begin     s = 4'b1101;    co = 2'b01;    end
        else if(    a == 4'b1111 && b == 4'b1101 && ci == 1'b1 )begin     s = 4'b1110;    co = 2'b01;    end
        else if(    a == 4'b1111 && b == 4'b1110 && ci == 1'b0 )begin     s = 4'b1110;    co = 2'b01;    end
        else if(    a == 4'b1111 && b == 4'b1110 && ci == 1'b1 )begin     s = 4'b0000;    co = 2'b10;    end
        else if(    a == 4'b1111 && b == 4'b1111 && ci == 1'b0 )begin     s = 4'b0000;    co = 2'b10;    end
        else if(    a == 4'b1111 && b == 4'b1111 && ci == 1'b1 )begin     s = 4'b0001;    co = 2'b10;    end
    end
endmodule