module xor_gate (A,B,C);
    input A,B;
    output C;
    
    xor(C,A,B);
    
endmodule