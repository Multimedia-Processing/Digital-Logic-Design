
`timescale 1ns/1ps

module T;
    reg Clk10M = 1'b0;
    reg Clr = 1'b1;
    reg Up = 1'b0;
    reg Down = 1'b0;
    wire Clk_o;
    wire [2:0] State;
    wire [14:0] Cnt;

    parameter PERIOD = 200;
    parameter real DUTY_CYCLE = 0.5;
    parameter OFFSET = 0;

    initial    // Clock process for Clk10M
    begin
        #OFFSET;
        forever
        begin
            Clk10M = 1'b0;
            #(PERIOD-(PERIOD*DUTY_CYCLE)) Clk10M = 1'b1;
            #(PERIOD*DUTY_CYCLE);
        end
    end

    buzzer UUT (
        .Clk10M(Clk10M),
        .Clr(Clr),
        .Up(Up),
        .Down(Down),
        .Clk_o(Clk_o),
        .State(State),
        .Cnt(Cnt));

    initial
    begin
      #56200 // Final time:  56200 ns
        $stop;
    end

    initial begin
        // -------------  Current Time:  285ns
        #285;
        Clr = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  2485ns
        #2200;
        Up = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  3485ns
        #1000;
        Up = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  5885ns
        #2400;
        Up = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  6885ns
        #1000;
        Up = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  9285ns
        #2400;
        Up = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  10285ns
        #1000;
        Up = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  12685ns
        #2400;
        Up = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  13685ns
        #1000;
        Up = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  16085ns
        #2400;
        Up = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  17085ns
        #1000;
        Up = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  19485ns
        #2400;
        Up = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  20485ns
        #1000;
        Up = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  22885ns
        #2400;
        Up = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  23885ns
        #1000;
        Up = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  27285ns
        #3400;
        Up = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  28685ns
        #1400;
        Down = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  29685ns
        #1000;
        Down = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  30685ns
        #1000;
        Up = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  32085ns
        #1400;
        Down = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  33085ns
        #1000;
        Down = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  34085ns
        #1000;
        Up = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  35485ns
        #1400;
        Down = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  36485ns
        #1000;
        Down = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  37485ns
        #1000;
        Up = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  38885ns
        #1400;
        Down = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  39885ns
        #1000;
        Down = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  42285ns
        #2400;
        Down = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  43285ns
        #1000;
        Down = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  44285ns
        #1000;
        Up = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  45685ns
        #1400;
        Down = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  46685ns
        #1000;
        Down = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  47685ns
        #1000;
        Up = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  49085ns
        #1400;
        Down = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  50085ns
        #1000;
        Down = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  51085ns
        #1000;
        Up = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  52285ns
        #1200;
        Up = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  53485ns
        #1200;
        Up = 1'b0;
        // -------------------------------------
    end

endmodule

