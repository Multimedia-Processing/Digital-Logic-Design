module NOR_GATE (c, a, b);

input a, b;
output c;

    nor(c, a, b);

endmodule