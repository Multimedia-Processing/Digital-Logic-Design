module NOT_GATE_A (c, a);

input a;
output c;

    not(c, a);

endmodule