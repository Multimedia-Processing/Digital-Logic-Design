module adder_4bit_case(a, b, ci, s, co);
    input [3:0] a,b;
    input ci;
    output [3:0] s;
    output [1:0] co;
    reg [3:0] s;
    reg [1:0] co;

    always@(a or b or ci)begin
        case({a, b, ci})
        //  a=0, b=0~F, c=0~1, truth table check ( OK )
        { 4'b0000 , 4'b0000 , 1'b0 }: begin     s = 4'b0000;    co = 2'b00;    end
        { 4'b0000 , 4'b0000 , 1'b1 }: begin     s = 4'b0001;    co = 2'b00;    end
        { 4'b0000 , 4'b0001 , 1'b0 }: begin     s = 4'b0001;    co = 2'b00;    end
        { 4'b0000 , 4'b0001 , 1'b1 }: begin     s = 4'b0010;    co = 2'b00;    end
        { 4'b0000 , 4'b0010 , 1'b0 }: begin     s = 4'b0010;    co = 2'b00;    end
        { 4'b0000 , 4'b0010 , 1'b1 }: begin     s = 4'b0011;    co = 2'b00;    end
        { 4'b0000 , 4'b0011 , 1'b0 }: begin     s = 4'b0011;    co = 2'b00;    end
        { 4'b0000 , 4'b0011 , 1'b1 }: begin     s = 4'b0100;    co = 2'b00;    end
        { 4'b0000 , 4'b0100 , 1'b0 }: begin     s = 4'b0100;    co = 2'b00;    end
        { 4'b0000 , 4'b0100 , 1'b1 }: begin     s = 4'b0101;    co = 2'b00;    end
        { 4'b0000 , 4'b0101 , 1'b0 }: begin     s = 4'b0101;    co = 2'b00;    end
        { 4'b0000 , 4'b0101 , 1'b1 }: begin     s = 4'b0110;    co = 2'b00;    end
        { 4'b0000 , 4'b0110 , 1'b0 }: begin     s = 4'b0110;    co = 2'b00;    end
        { 4'b0000 , 4'b0110 , 1'b1 }: begin     s = 4'b0111;    co = 2'b00;    end
        { 4'b0000 , 4'b0111 , 1'b0 }: begin     s = 4'b0111;    co = 2'b00;    end
        { 4'b0000 , 4'b0111 , 1'b1 }: begin     s = 4'b1000;    co = 2'b00;    end
        { 4'b0000 , 4'b1000 , 1'b0 }: begin     s = 4'b1000;    co = 2'b00;    end
        { 4'b0000 , 4'b1000 , 1'b1 }: begin     s = 4'b1001;    co = 2'b00;    end
        { 4'b0000 , 4'b1001 , 1'b0 }: begin     s = 4'b1001;    co = 2'b00;    end
        { 4'b0000 , 4'b1001 , 1'b1 }: begin     s = 4'b1010;    co = 2'b00;    end
        { 4'b0000 , 4'b1010 , 1'b0 }: begin     s = 4'b1010;    co = 2'b00;    end
        { 4'b0000 , 4'b1010 , 1'b1 }: begin     s = 4'b1011;    co = 2'b00;    end
        { 4'b0000 , 4'b1011 , 1'b0 }: begin     s = 4'b1011;    co = 2'b00;    end
        { 4'b0000 , 4'b1011 , 1'b1 }: begin     s = 4'b1100;    co = 2'b00;    end
        { 4'b0000 , 4'b1100 , 1'b0 }: begin     s = 4'b1100;    co = 2'b00;    end
        { 4'b0000 , 4'b1100 , 1'b1 }: begin     s = 4'b1101;    co = 2'b00;    end
        { 4'b0000 , 4'b1101 , 1'b0 }: begin     s = 4'b1101;    co = 2'b00;    end
        { 4'b0000 , 4'b1101 , 1'b1 }: begin     s = 4'b1110;    co = 2'b00;    end
        { 4'b0000 , 4'b1110 , 1'b0 }: begin     s = 4'b1110;    co = 2'b00;    end
        { 4'b0000 , 4'b1110 , 1'b1 }: begin     s = 4'b1111;    co = 2'b00;    end
        { 4'b0000 , 4'b1111 , 1'b0 }: begin     s = 4'b1111;    co = 2'b00;    end
        { 4'b0000 , 4'b1111 , 1'b1 }: begin     s = 4'b0000;    co = 2'b01;    end
        //  a=1, b=0~F, c=0~1, truth table check ( OK )
        { 4'b0001 , 4'b0000 , 1'b0 }: begin     s = 4'b0001;    co = 2'b00;    end
        { 4'b0001 , 4'b0000 , 1'b1 }: begin     s = 4'b0010;    co = 2'b00;    end
        { 4'b0001 , 4'b0001 , 1'b0 }: begin     s = 4'b0010;    co = 2'b00;    end
        { 4'b0001 , 4'b0001 , 1'b1 }: begin     s = 4'b0011;    co = 2'b00;    end
        { 4'b0001 , 4'b0010 , 1'b0 }: begin     s = 4'b0011;    co = 2'b00;    end
        { 4'b0001 , 4'b0010 , 1'b1 }: begin     s = 4'b0100;    co = 2'b00;    end
        { 4'b0001 , 4'b0011 , 1'b0 }: begin     s = 4'b0100;    co = 2'b00;    end
        { 4'b0001 , 4'b0011 , 1'b1 }: begin     s = 4'b0101;    co = 2'b00;    end
        { 4'b0001 , 4'b0100 , 1'b0 }: begin     s = 4'b0101;    co = 2'b00;    end
        { 4'b0001 , 4'b0100 , 1'b1 }: begin     s = 4'b0110;    co = 2'b00;    end
        { 4'b0001 , 4'b0101 , 1'b0 }: begin     s = 4'b0110;    co = 2'b00;    end
        { 4'b0001 , 4'b0101 , 1'b1 }: begin     s = 4'b0111;    co = 2'b00;    end
        { 4'b0001 , 4'b0110 , 1'b0 }: begin     s = 4'b0111;    co = 2'b00;    end
        { 4'b0001 , 4'b0110 , 1'b1 }: begin     s = 4'b1000;    co = 2'b00;    end
        { 4'b0001 , 4'b0111 , 1'b0 }: begin     s = 4'b1000;    co = 2'b00;    end
        { 4'b0001 , 4'b0111 , 1'b1 }: begin     s = 4'b1001;    co = 2'b00;    end
        { 4'b0001 , 4'b1000 , 1'b0 }: begin     s = 4'b1001;    co = 2'b00;    end
        { 4'b0001 , 4'b1000 , 1'b1 }: begin     s = 4'b1010;    co = 2'b00;    end
        { 4'b0001 , 4'b1001 , 1'b0 }: begin     s = 4'b1010;    co = 2'b00;    end
        { 4'b0001 , 4'b1001 , 1'b1 }: begin     s = 4'b1011;    co = 2'b00;    end
        { 4'b0001 , 4'b1010 , 1'b0 }: begin     s = 4'b1011;    co = 2'b00;    end
        { 4'b0001 , 4'b1010 , 1'b1 }: begin     s = 4'b1100;    co = 2'b00;    end
        { 4'b0001 , 4'b1011 , 1'b0 }: begin     s = 4'b1100;    co = 2'b00;    end
        { 4'b0001 , 4'b1011 , 1'b1 }: begin     s = 4'b1101;    co = 2'b00;    end
        { 4'b0001 , 4'b1100 , 1'b0 }: begin     s = 4'b1101;    co = 2'b00;    end
        { 4'b0001 , 4'b1100 , 1'b1 }: begin     s = 4'b1110;    co = 2'b00;    end
        { 4'b0001 , 4'b1101 , 1'b0 }: begin     s = 4'b1110;    co = 2'b00;    end
        { 4'b0001 , 4'b1101 , 1'b1 }: begin     s = 4'b1111;    co = 2'b00;    end
        { 4'b0001 , 4'b1110 , 1'b0 }: begin     s = 4'b1111;    co = 2'b00;    end
        { 4'b0001 , 4'b1110 , 1'b1 }: begin     s = 4'b0000;    co = 2'b01;    end
        { 4'b0001 , 4'b1111 , 1'b0 }: begin     s = 4'b0000;    co = 2'b01;    end
        { 4'b0001 , 4'b1111 , 1'b1 }: begin     s = 4'b0001;    co = 2'b01;    end
        //  a=2, b=0~F, c=0~1, truth table check ( OK )
        { 4'b0010 , 4'b0000 , 1'b0 }: begin     s = 4'b0010;    co = 2'b00;    end
        { 4'b0010 , 4'b0000 , 1'b1 }: begin     s = 4'b0011;    co = 2'b00;    end
        { 4'b0010 , 4'b0001 , 1'b0 }: begin     s = 4'b0011;    co = 2'b00;    end
        { 4'b0010 , 4'b0001 , 1'b1 }: begin     s = 4'b0100;    co = 2'b00;    end
        { 4'b0010 , 4'b0010 , 1'b0 }: begin     s = 4'b0100;    co = 2'b00;    end
        { 4'b0010 , 4'b0010 , 1'b1 }: begin     s = 4'b0101;    co = 2'b00;    end
        { 4'b0010 , 4'b0011 , 1'b0 }: begin     s = 4'b0101;    co = 2'b00;    end
        { 4'b0010 , 4'b0011 , 1'b1 }: begin     s = 4'b0110;    co = 2'b00;    end
        { 4'b0010 , 4'b0100 , 1'b0 }: begin     s = 4'b0110;    co = 2'b00;    end
        { 4'b0010 , 4'b0100 , 1'b1 }: begin     s = 4'b0111;    co = 2'b00;    end
        { 4'b0010 , 4'b0101 , 1'b0 }: begin     s = 4'b0111;    co = 2'b00;    end
        { 4'b0010 , 4'b0101 , 1'b1 }: begin     s = 4'b1000;    co = 2'b00;    end
        { 4'b0010 , 4'b0110 , 1'b0 }: begin     s = 4'b1000;    co = 2'b00;    end
        { 4'b0010 , 4'b0110 , 1'b1 }: begin     s = 4'b1001;    co = 2'b00;    end
        { 4'b0010 , 4'b0111 , 1'b0 }: begin     s = 4'b1001;    co = 2'b00;    end
        { 4'b0010 , 4'b0111 , 1'b1 }: begin     s = 4'b1010;    co = 2'b00;    end
        { 4'b0010 , 4'b1000 , 1'b0 }: begin     s = 4'b1010;    co = 2'b00;    end
        { 4'b0010 , 4'b1000 , 1'b1 }: begin     s = 4'b1011;    co = 2'b00;    end
        { 4'b0010 , 4'b1001 , 1'b0 }: begin     s = 4'b1011;    co = 2'b00;    end
        { 4'b0010 , 4'b1001 , 1'b1 }: begin     s = 4'b1100;    co = 2'b00;    end
        { 4'b0010 , 4'b1010 , 1'b0 }: begin     s = 4'b1100;    co = 2'b00;    end
        { 4'b0010 , 4'b1010 , 1'b1 }: begin     s = 4'b1101;    co = 2'b00;    end
        { 4'b0010 , 4'b1011 , 1'b0 }: begin     s = 4'b1101;    co = 2'b00;    end
        { 4'b0010 , 4'b1011 , 1'b1 }: begin     s = 4'b1110;    co = 2'b00;    end
        { 4'b0010 , 4'b1100 , 1'b0 }: begin     s = 4'b1110;    co = 2'b00;    end
        { 4'b0010 , 4'b1100 , 1'b1 }: begin     s = 4'b1111;    co = 2'b00;    end
        { 4'b0010 , 4'b1101 , 1'b0 }: begin     s = 4'b1111;    co = 2'b00;    end
        { 4'b0010 , 4'b1101 , 1'b1 }: begin     s = 4'b0000;    co = 2'b01;    end
        { 4'b0010 , 4'b1110 , 1'b0 }: begin     s = 4'b0000;    co = 2'b01;    end
        { 4'b0010 , 4'b1110 , 1'b1 }: begin     s = 4'b0001;    co = 2'b01;    end
        { 4'b0010 , 4'b1111 , 1'b0 }: begin     s = 4'b0001;    co = 2'b01;    end
        { 4'b0010 , 4'b1111 , 1'b1 }: begin     s = 4'b0010;    co = 2'b01;    end
        //  a=3, b=0~F, c=0~1, truth table check ( OK )
        { 4'b0011 , 4'b0000 , 1'b0 }: begin     s = 4'b0011;    co = 2'b00;    end
        { 4'b0011 , 4'b0000 , 1'b1 }: begin     s = 4'b0100;    co = 2'b00;    end
        { 4'b0011 , 4'b0001 , 1'b0 }: begin     s = 4'b0100;    co = 2'b00;    end
        { 4'b0011 , 4'b0001 , 1'b1 }: begin     s = 4'b0101;    co = 2'b00;    end
        { 4'b0011 , 4'b0010 , 1'b0 }: begin     s = 4'b0101;    co = 2'b00;    end
        { 4'b0011 , 4'b0010 , 1'b1 }: begin     s = 4'b0110;    co = 2'b00;    end
        { 4'b0011 , 4'b0011 , 1'b0 }: begin     s = 4'b0110;    co = 2'b00;    end
        { 4'b0011 , 4'b0011 , 1'b1 }: begin     s = 4'b0111;    co = 2'b00;    end
        { 4'b0011 , 4'b0100 , 1'b0 }: begin     s = 4'b0111;    co = 2'b00;    end
        { 4'b0011 , 4'b0100 , 1'b1 }: begin     s = 4'b1000;    co = 2'b00;    end
        { 4'b0011 , 4'b0101 , 1'b0 }: begin     s = 4'b1000;    co = 2'b00;    end
        { 4'b0011 , 4'b0101 , 1'b1 }: begin     s = 4'b1001;    co = 2'b00;    end
        { 4'b0011 , 4'b0110 , 1'b0 }: begin     s = 4'b1001;    co = 2'b00;    end
        { 4'b0011 , 4'b0110 , 1'b1 }: begin     s = 4'b1010;    co = 2'b00;    end
        { 4'b0011 , 4'b0111 , 1'b0 }: begin     s = 4'b1010;    co = 2'b00;    end
        { 4'b0011 , 4'b0111 , 1'b1 }: begin     s = 4'b1011;    co = 2'b00;    end
        { 4'b0011 , 4'b1000 , 1'b0 }: begin     s = 4'b1011;    co = 2'b00;    end
        { 4'b0011 , 4'b1000 , 1'b1 }: begin     s = 4'b1100;    co = 2'b00;    end
        { 4'b0011 , 4'b1001 , 1'b0 }: begin     s = 4'b1100;    co = 2'b00;    end
        { 4'b0011 , 4'b1001 , 1'b1 }: begin     s = 4'b1101;    co = 2'b00;    end
        { 4'b0011 , 4'b1010 , 1'b0 }: begin     s = 4'b1101;    co = 2'b00;    end
        { 4'b0011 , 4'b1010 , 1'b1 }: begin     s = 4'b1110;    co = 2'b00;    end
        { 4'b0011 , 4'b1011 , 1'b0 }: begin     s = 4'b1110;    co = 2'b00;    end
        { 4'b0011 , 4'b1011 , 1'b1 }: begin     s = 4'b1111;    co = 2'b00;    end
        { 4'b0011 , 4'b1100 , 1'b0 }: begin     s = 4'b1111;    co = 2'b00;    end
        { 4'b0011 , 4'b1100 , 1'b1 }: begin     s = 4'b0000;    co = 2'b01;    end
        { 4'b0011 , 4'b1101 , 1'b0 }: begin     s = 4'b0000;    co = 2'b01;    end
        { 4'b0011 , 4'b1101 , 1'b1 }: begin     s = 4'b0011;    co = 2'b01;    end
        { 4'b0011 , 4'b1110 , 1'b0 }: begin     s = 4'b0011;    co = 2'b01;    end
        { 4'b0011 , 4'b1110 , 1'b1 }: begin     s = 4'b0010;    co = 2'b01;    end
        { 4'b0011 , 4'b1111 , 1'b0 }: begin     s = 4'b0010;    co = 2'b01;    end
        { 4'b0011 , 4'b1111 , 1'b1 }: begin     s = 4'b0011;    co = 2'b01;    end
        //  a=4, b=0~F, c=0~1, truth table check ( OK )
        { 4'b0100 , 4'b0000 , 1'b0 }: begin     s = 4'b0100;    co = 2'b00;    end
        { 4'b0100 , 4'b0000 , 1'b1 }: begin     s = 4'b0101;    co = 2'b00;    end
        { 4'b0100 , 4'b0001 , 1'b0 }: begin     s = 4'b0101;    co = 2'b00;    end
        { 4'b0100 , 4'b0001 , 1'b1 }: begin     s = 4'b0110;    co = 2'b00;    end
        { 4'b0100 , 4'b0010 , 1'b0 }: begin     s = 4'b0110;    co = 2'b00;    end
        { 4'b0100 , 4'b0010 , 1'b1 }: begin     s = 4'b0111;    co = 2'b00;    end
        { 4'b0100 , 4'b0011 , 1'b0 }: begin     s = 4'b0111;    co = 2'b00;    end
        { 4'b0100 , 4'b0011 , 1'b1 }: begin     s = 4'b1000;    co = 2'b00;    end
        { 4'b0100 , 4'b0100 , 1'b0 }: begin     s = 4'b1000;    co = 2'b00;    end
        { 4'b0100 , 4'b0100 , 1'b1 }: begin     s = 4'b1001;    co = 2'b00;    end
        { 4'b0100 , 4'b0101 , 1'b0 }: begin     s = 4'b1001;    co = 2'b00;    end
        { 4'b0100 , 4'b0101 , 1'b1 }: begin     s = 4'b1010;    co = 2'b00;    end
        { 4'b0100 , 4'b0110 , 1'b0 }: begin     s = 4'b1010;    co = 2'b00;    end
        { 4'b0100 , 4'b0110 , 1'b1 }: begin     s = 4'b1011;    co = 2'b00;    end
        { 4'b0100 , 4'b0111 , 1'b0 }: begin     s = 4'b1011;    co = 2'b00;    end
        { 4'b0100 , 4'b0111 , 1'b1 }: begin     s = 4'b1100;    co = 2'b00;    end
        { 4'b0100 , 4'b1000 , 1'b0 }: begin     s = 4'b1100;    co = 2'b00;    end
        { 4'b0100 , 4'b1000 , 1'b1 }: begin     s = 4'b1101;    co = 2'b00;    end
        { 4'b0100 , 4'b1001 , 1'b0 }: begin     s = 4'b1101;    co = 2'b00;    end
        { 4'b0100 , 4'b1001 , 1'b1 }: begin     s = 4'b1110;    co = 2'b00;    end
        { 4'b0100 , 4'b1010 , 1'b0 }: begin     s = 4'b1110;    co = 2'b00;    end
        { 4'b0100 , 4'b1010 , 1'b1 }: begin     s = 4'b1111;    co = 2'b00;    end
        { 4'b0100 , 4'b1011 , 1'b0 }: begin     s = 4'b1111;    co = 2'b00;    end
        { 4'b0100 , 4'b1011 , 1'b1 }: begin     s = 4'b0000;    co = 2'b01;    end
        { 4'b0100 , 4'b1100 , 1'b0 }: begin     s = 4'b0000;    co = 2'b01;    end
        { 4'b0100 , 4'b1100 , 1'b1 }: begin     s = 4'b0001;    co = 2'b01;    end
        { 4'b0100 , 4'b1101 , 1'b0 }: begin     s = 4'b0001;    co = 2'b01;    end
        { 4'b0100 , 4'b1101 , 1'b1 }: begin     s = 4'b0010;    co = 2'b01;    end
        { 4'b0100 , 4'b1110 , 1'b0 }: begin     s = 4'b0010;    co = 2'b01;    end
        { 4'b0100 , 4'b1110 , 1'b1 }: begin     s = 4'b0011;    co = 2'b01;    end
        { 4'b0100 , 4'b1111 , 1'b0 }: begin     s = 4'b0011;    co = 2'b01;    end
        { 4'b0100 , 4'b1111 , 1'b1 }: begin     s = 4'b0100;    co = 2'b01;    end
        //  a=5, b=0~F, c=0~1, truth table check ( OK )
        { 4'b0101 , 4'b0000 , 1'b0 }: begin     s = 4'b0101;    co = 2'b00;    end
        { 4'b0101 , 4'b0000 , 1'b1 }: begin     s = 4'b0110;    co = 2'b00;    end
        { 4'b0101 , 4'b0001 , 1'b0 }: begin     s = 4'b0110;    co = 2'b00;    end
        { 4'b0101 , 4'b0001 , 1'b1 }: begin     s = 4'b0111;    co = 2'b00;    end
        { 4'b0101 , 4'b0010 , 1'b0 }: begin     s = 4'b0111;    co = 2'b00;    end
        { 4'b0101 , 4'b0010 , 1'b1 }: begin     s = 4'b1000;    co = 2'b00;    end
        { 4'b0101 , 4'b0011 , 1'b0 }: begin     s = 4'b1000;    co = 2'b00;    end
        { 4'b0101 , 4'b0011 , 1'b1 }: begin     s = 4'b1001;    co = 2'b00;    end
        { 4'b0101 , 4'b0100 , 1'b0 }: begin     s = 4'b1001;    co = 2'b00;    end
        { 4'b0101 , 4'b0100 , 1'b1 }: begin     s = 4'b1010;    co = 2'b00;    end
        { 4'b0101 , 4'b0101 , 1'b0 }: begin     s = 4'b1010;    co = 2'b00;    end
        { 4'b0101 , 4'b0101 , 1'b1 }: begin     s = 4'b1011;    co = 2'b00;    end
        { 4'b0101 , 4'b0110 , 1'b0 }: begin     s = 4'b1011;    co = 2'b00;    end
        { 4'b0101 , 4'b0110 , 1'b1 }: begin     s = 4'b1100;    co = 2'b00;    end
        { 4'b0101 , 4'b0111 , 1'b0 }: begin     s = 4'b1100;    co = 2'b00;    end
        { 4'b0101 , 4'b0111 , 1'b1 }: begin     s = 4'b1101;    co = 2'b00;    end
        { 4'b0101 , 4'b1000 , 1'b0 }: begin     s = 4'b1101;    co = 2'b00;    end
        { 4'b0101 , 4'b1000 , 1'b1 }: begin     s = 4'b1110;    co = 2'b00;    end
        { 4'b0101 , 4'b1001 , 1'b0 }: begin     s = 4'b1110;    co = 2'b00;    end
        { 4'b0101 , 4'b1001 , 1'b1 }: begin     s = 4'b1111;    co = 2'b00;    end
        { 4'b0101 , 4'b1010 , 1'b0 }: begin     s = 4'b1111;    co = 2'b00;    end
        { 4'b0101 , 4'b1010 , 1'b1 }: begin     s = 4'b0000;    co = 2'b01;    end
        { 4'b0101 , 4'b1011 , 1'b0 }: begin     s = 4'b0000;    co = 2'b01;    end
        { 4'b0101 , 4'b1011 , 1'b1 }: begin     s = 4'b0001;    co = 2'b01;    end
        { 4'b0101 , 4'b1100 , 1'b0 }: begin     s = 4'b0001;    co = 2'b01;    end
        { 4'b0101 , 4'b1100 , 1'b1 }: begin     s = 4'b0010;    co = 2'b01;    end
        { 4'b0101 , 4'b1101 , 1'b0 }: begin     s = 4'b0010;    co = 2'b01;    end
        { 4'b0101 , 4'b1101 , 1'b1 }: begin     s = 4'b0011;    co = 2'b01;    end
        { 4'b0101 , 4'b1110 , 1'b0 }: begin     s = 4'b0011;    co = 2'b01;    end
        { 4'b0101 , 4'b1110 , 1'b1 }: begin     s = 4'b0100;    co = 2'b01;    end
        { 4'b0101 , 4'b1111 , 1'b0 }: begin     s = 4'b0100;    co = 2'b01;    end
        { 4'b0101 , 4'b1111 , 1'b1 }: begin     s = 4'b0101;    co = 2'b01;    end
        //  a=6, b=0~F, c=0~1, truth table check ( OK )
        { 4'b0110 , 4'b0000 , 1'b0 }: begin     s = 4'b0110;    co = 2'b00;    end
        { 4'b0110 , 4'b0000 , 1'b1 }: begin     s = 4'b0111;    co = 2'b00;    end
        { 4'b0110 , 4'b0001 , 1'b0 }: begin     s = 4'b0111;    co = 2'b00;    end
        { 4'b0110 , 4'b0001 , 1'b1 }: begin     s = 4'b1000;    co = 2'b00;    end
        { 4'b0110 , 4'b0010 , 1'b0 }: begin     s = 4'b1000;    co = 2'b00;    end
        { 4'b0110 , 4'b0010 , 1'b1 }: begin     s = 4'b1001;    co = 2'b00;    end
        { 4'b0110 , 4'b0011 , 1'b0 }: begin     s = 4'b1001;    co = 2'b00;    end
        { 4'b0110 , 4'b0011 , 1'b1 }: begin     s = 4'b1010;    co = 2'b00;    end
        { 4'b0110 , 4'b0100 , 1'b0 }: begin     s = 4'b1010;    co = 2'b00;    end
        { 4'b0110 , 4'b0100 , 1'b1 }: begin     s = 4'b1011;    co = 2'b00;    end
        { 4'b0110 , 4'b0101 , 1'b0 }: begin     s = 4'b1011;    co = 2'b00;    end
        { 4'b0110 , 4'b0101 , 1'b1 }: begin     s = 4'b1100;    co = 2'b00;    end
        { 4'b0110 , 4'b0110 , 1'b0 }: begin     s = 4'b1100;    co = 2'b00;    end
        { 4'b0110 , 4'b0110 , 1'b1 }: begin     s = 4'b1101;    co = 2'b00;    end
        { 4'b0110 , 4'b0111 , 1'b0 }: begin     s = 4'b1101;    co = 2'b00;    end
        { 4'b0110 , 4'b0111 , 1'b1 }: begin     s = 4'b1110;    co = 2'b00;    end
        { 4'b0110 , 4'b1000 , 1'b0 }: begin     s = 4'b1110;    co = 2'b00;    end
        { 4'b0110 , 4'b1000 , 1'b1 }: begin     s = 4'b1111;    co = 2'b00;    end
        { 4'b0110 , 4'b1001 , 1'b0 }: begin     s = 4'b1111;    co = 2'b00;    end
        { 4'b0110 , 4'b1001 , 1'b1 }: begin     s = 4'b0000;    co = 2'b01;    end
        { 4'b0110 , 4'b1010 , 1'b0 }: begin     s = 4'b0000;    co = 2'b01;    end
        { 4'b0110 , 4'b1010 , 1'b1 }: begin     s = 4'b0001;    co = 2'b01;    end
        { 4'b0110 , 4'b1011 , 1'b0 }: begin     s = 4'b0001;    co = 2'b01;    end
        { 4'b0110 , 4'b1011 , 1'b1 }: begin     s = 4'b0010;    co = 2'b01;    end
        { 4'b0110 , 4'b1100 , 1'b0 }: begin     s = 4'b0010;    co = 2'b01;    end
        { 4'b0110 , 4'b1100 , 1'b1 }: begin     s = 4'b0011;    co = 2'b01;    end
        { 4'b0110 , 4'b1101 , 1'b0 }: begin     s = 4'b0011;    co = 2'b01;    end
        { 4'b0110 , 4'b1101 , 1'b1 }: begin     s = 4'b0100;    co = 2'b01;    end
        { 4'b0110 , 4'b1110 , 1'b0 }: begin     s = 4'b0100;    co = 2'b01;    end
        { 4'b0110 , 4'b1110 , 1'b1 }: begin     s = 4'b0101;    co = 2'b01;    end
        { 4'b0110 , 4'b1111 , 1'b0 }: begin     s = 4'b0101;    co = 2'b01;    end
        { 4'b0110 , 4'b1111 , 1'b1 }: begin     s = 4'b0110;    co = 2'b01;    end
        //  a=7, b=0~F, c=0~1, truth table check ( OK )
        { 4'b0111 , 4'b0000 , 1'b0 }: begin     s = 4'b0111;    co = 2'b00;    end
        { 4'b0111 , 4'b0000 , 1'b1 }: begin     s = 4'b1000;    co = 2'b00;    end
        { 4'b0111 , 4'b0001 , 1'b0 }: begin     s = 4'b1000;    co = 2'b00;    end
        { 4'b0111 , 4'b0001 , 1'b1 }: begin     s = 4'b1001;    co = 2'b00;    end
        { 4'b0111 , 4'b0010 , 1'b0 }: begin     s = 4'b1001;    co = 2'b00;    end
        { 4'b0111 , 4'b0010 , 1'b1 }: begin     s = 4'b1010;    co = 2'b00;    end
        { 4'b0111 , 4'b0011 , 1'b0 }: begin     s = 4'b1010;    co = 2'b00;    end
        { 4'b0111 , 4'b0011 , 1'b1 }: begin     s = 4'b1011;    co = 2'b00;    end
        { 4'b0111 , 4'b0100 , 1'b0 }: begin     s = 4'b1011;    co = 2'b00;    end
        { 4'b0111 , 4'b0100 , 1'b1 }: begin     s = 4'b1100;    co = 2'b00;    end
        { 4'b0111 , 4'b0101 , 1'b0 }: begin     s = 4'b1100;    co = 2'b00;    end
        { 4'b0111 , 4'b0101 , 1'b1 }: begin     s = 4'b1101;    co = 2'b00;    end
        { 4'b0111 , 4'b0110 , 1'b0 }: begin     s = 4'b1101;    co = 2'b00;    end
        { 4'b0111 , 4'b0110 , 1'b1 }: begin     s = 4'b1110;    co = 2'b00;    end
        { 4'b0111 , 4'b0111 , 1'b0 }: begin     s = 4'b1110;    co = 2'b00;    end
        { 4'b0111 , 4'b0111 , 1'b1 }: begin     s = 4'b1111;    co = 2'b00;    end
        { 4'b0111 , 4'b1000 , 1'b0 }: begin     s = 4'b1111;    co = 2'b00;    end
        { 4'b0111 , 4'b1000 , 1'b1 }: begin     s = 4'b0000;    co = 2'b01;    end
        { 4'b0111 , 4'b1001 , 1'b0 }: begin     s = 4'b0000;    co = 2'b01;    end
        { 4'b0111 , 4'b1001 , 1'b1 }: begin     s = 4'b0001;    co = 2'b01;    end
        { 4'b0111 , 4'b1010 , 1'b0 }: begin     s = 4'b0001;    co = 2'b01;    end
        { 4'b0111 , 4'b1010 , 1'b1 }: begin     s = 4'b0010;    co = 2'b01;    end
        { 4'b0111 , 4'b1011 , 1'b0 }: begin     s = 4'b0010;    co = 2'b01;    end
        { 4'b0111 , 4'b1011 , 1'b1 }: begin     s = 4'b0011;    co = 2'b01;    end
        { 4'b0111 , 4'b1100 , 1'b0 }: begin     s = 4'b0011;    co = 2'b01;    end
        { 4'b0111 , 4'b1100 , 1'b1 }: begin     s = 4'b0100;    co = 2'b01;    end
        { 4'b0111 , 4'b1101 , 1'b0 }: begin     s = 4'b0100;    co = 2'b01;    end
        { 4'b0111 , 4'b1101 , 1'b1 }: begin     s = 4'b0101;    co = 2'b01;    end
        { 4'b0111 , 4'b1110 , 1'b0 }: begin     s = 4'b0101;    co = 2'b01;    end
        { 4'b0111 , 4'b1110 , 1'b1 }: begin     s = 4'b0110;    co = 2'b01;    end
        { 4'b0111 , 4'b1111 , 1'b0 }: begin     s = 4'b0110;    co = 2'b01;    end
        { 4'b0111 , 4'b1111 , 1'b1 }: begin     s = 4'b0111;    co = 2'b01;    end
        //  a=8, b=0~F, c=0~1, truth table check ( OK )
        { 4'b1000 , 4'b0000 , 1'b0 }: begin     s = 4'b1000;    co = 2'b00;    end
        { 4'b1000 , 4'b0000 , 1'b1 }: begin     s = 4'b1001;    co = 2'b00;    end
        { 4'b1000 , 4'b0001 , 1'b0 }: begin     s = 4'b1001;    co = 2'b00;    end
        { 4'b1000 , 4'b0001 , 1'b1 }: begin     s = 4'b1010;    co = 2'b00;    end
        { 4'b1000 , 4'b0010 , 1'b0 }: begin     s = 4'b1010;    co = 2'b00;    end
        { 4'b1000 , 4'b0010 , 1'b1 }: begin     s = 4'b1011;    co = 2'b00;    end
        { 4'b1000 , 4'b0011 , 1'b0 }: begin     s = 4'b1011;    co = 2'b00;    end
        { 4'b1000 , 4'b0011 , 1'b1 }: begin     s = 4'b1100;    co = 2'b00;    end
        { 4'b1000 , 4'b0100 , 1'b0 }: begin     s = 4'b1100;    co = 2'b00;    end
        { 4'b1000 , 4'b0100 , 1'b1 }: begin     s = 4'b1101;    co = 2'b00;    end
        { 4'b1000 , 4'b0101 , 1'b0 }: begin     s = 4'b1101;    co = 2'b00;    end
        { 4'b1000 , 4'b0101 , 1'b1 }: begin     s = 4'b1110;    co = 2'b00;    end
        { 4'b1000 , 4'b0110 , 1'b0 }: begin     s = 4'b1110;    co = 2'b00;    end
        { 4'b1000 , 4'b0110 , 1'b1 }: begin     s = 4'b1111;    co = 2'b00;    end
        { 4'b1000 , 4'b0111 , 1'b0 }: begin     s = 4'b1111;    co = 2'b00;    end
        { 4'b1000 , 4'b0111 , 1'b1 }: begin     s = 4'b0000;    co = 2'b01;    end
        { 4'b1000 , 4'b1000 , 1'b0 }: begin     s = 4'b0000;    co = 2'b01;    end
        { 4'b1000 , 4'b1000 , 1'b1 }: begin     s = 4'b0001;    co = 2'b01;    end
        { 4'b1000 , 4'b1001 , 1'b0 }: begin     s = 4'b0001;    co = 2'b01;    end
        { 4'b1000 , 4'b1001 , 1'b1 }: begin     s = 4'b0010;    co = 2'b01;    end
        { 4'b1000 , 4'b1010 , 1'b0 }: begin     s = 4'b0010;    co = 2'b01;    end
        { 4'b1000 , 4'b1010 , 1'b1 }: begin     s = 4'b0011;    co = 2'b01;    end
        { 4'b1000 , 4'b1011 , 1'b0 }: begin     s = 4'b0011;    co = 2'b01;    end
        { 4'b1000 , 4'b1011 , 1'b1 }: begin     s = 4'b0100;    co = 2'b01;    end
        { 4'b1000 , 4'b1100 , 1'b0 }: begin     s = 4'b0100;    co = 2'b01;    end
        { 4'b1000 , 4'b1100 , 1'b1 }: begin     s = 4'b0101;    co = 2'b01;    end
        { 4'b1000 , 4'b1101 , 1'b0 }: begin     s = 4'b0101;    co = 2'b01;    end
        { 4'b1000 , 4'b1101 , 1'b1 }: begin     s = 4'b0110;    co = 2'b01;    end
        { 4'b1000 , 4'b1110 , 1'b0 }: begin     s = 4'b0110;    co = 2'b01;    end
        { 4'b1000 , 4'b1110 , 1'b1 }: begin     s = 4'b0111;    co = 2'b01;    end
        { 4'b1000 , 4'b1111 , 1'b0 }: begin     s = 4'b0111;    co = 2'b01;    end
        { 4'b1000 , 4'b1111 , 1'b1 }: begin     s = 4'b1000;    co = 2'b01;    end
        //  a=9, b=0~F, c=0~1, truth table check ( OK )
        { 4'b1001 , 4'b0000 , 1'b0 }: begin     s = 4'b1001;    co = 2'b00;    end
        { 4'b1001 , 4'b0000 , 1'b1 }: begin     s = 4'b1010;    co = 2'b00;    end
        { 4'b1001 , 4'b0001 , 1'b0 }: begin     s = 4'b1010;    co = 2'b00;    end
        { 4'b1001 , 4'b0001 , 1'b1 }: begin     s = 4'b1011;    co = 2'b00;    end
        { 4'b1001 , 4'b0010 , 1'b0 }: begin     s = 4'b1011;    co = 2'b00;    end
        { 4'b1001 , 4'b0010 , 1'b1 }: begin     s = 4'b1100;    co = 2'b00;    end
        { 4'b1001 , 4'b0011 , 1'b0 }: begin     s = 4'b1100;    co = 2'b00;    end
        { 4'b1001 , 4'b0011 , 1'b1 }: begin     s = 4'b1101;    co = 2'b00;    end
        { 4'b1001 , 4'b0100 , 1'b0 }: begin     s = 4'b1101;    co = 2'b00;    end
        { 4'b1001 , 4'b0100 , 1'b1 }: begin     s = 4'b1110;    co = 2'b00;    end
        { 4'b1001 , 4'b0101 , 1'b0 }: begin     s = 4'b1110;    co = 2'b00;    end
        { 4'b1001 , 4'b0101 , 1'b1 }: begin     s = 4'b1111;    co = 2'b00;    end
        { 4'b1001 , 4'b0110 , 1'b0 }: begin     s = 4'b1111;    co = 2'b00;    end
        { 4'b1001 , 4'b0110 , 1'b1 }: begin     s = 4'b0000;    co = 2'b01;    end
        { 4'b1001 , 4'b0111 , 1'b0 }: begin     s = 4'b0000;    co = 2'b01;    end
        { 4'b1001 , 4'b0111 , 1'b1 }: begin     s = 4'b0001;    co = 2'b01;    end
        { 4'b1001 , 4'b1000 , 1'b0 }: begin     s = 4'b0001;    co = 2'b01;    end
        { 4'b1001 , 4'b1000 , 1'b1 }: begin     s = 4'b0010;    co = 2'b01;    end
        { 4'b1001 , 4'b1001 , 1'b0 }: begin     s = 4'b0010;    co = 2'b01;    end
        { 4'b1001 , 4'b1001 , 1'b1 }: begin     s = 4'b0011;    co = 2'b01;    end
        { 4'b1001 , 4'b1010 , 1'b0 }: begin     s = 4'b0011;    co = 2'b01;    end
        { 4'b1001 , 4'b1010 , 1'b1 }: begin     s = 4'b0100;    co = 2'b01;    end
        { 4'b1001 , 4'b1011 , 1'b0 }: begin     s = 4'b0100;    co = 2'b01;    end
        { 4'b1001 , 4'b1011 , 1'b1 }: begin     s = 4'b0101;    co = 2'b01;    end
        { 4'b1001 , 4'b1100 , 1'b0 }: begin     s = 4'b0101;    co = 2'b01;    end
        { 4'b1001 , 4'b1100 , 1'b1 }: begin     s = 4'b0110;    co = 2'b01;    end
        { 4'b1001 , 4'b1101 , 1'b0 }: begin     s = 4'b0110;    co = 2'b01;    end
        { 4'b1001 , 4'b1101 , 1'b1 }: begin     s = 4'b0111;    co = 2'b01;    end
        { 4'b1001 , 4'b1110 , 1'b0 }: begin     s = 4'b0111;    co = 2'b01;    end
        { 4'b1001 , 4'b1110 , 1'b1 }: begin     s = 4'b1000;    co = 2'b01;    end
        { 4'b1001 , 4'b1111 , 1'b0 }: begin     s = 4'b1000;    co = 2'b01;    end
        { 4'b1001 , 4'b1111 , 1'b1 }: begin     s = 4'b1001;    co = 2'b01;    end
        //  a=A, b=0~F, c=0~1, truth table check ( OK )
        { 4'b1010 , 4'b0000 , 1'b0 }: begin     s = 4'b1010;    co = 2'b00;    end
        { 4'b1010 , 4'b0000 , 1'b1 }: begin     s = 4'b1011;    co = 2'b00;    end
        { 4'b1010 , 4'b0001 , 1'b0 }: begin     s = 4'b1011;    co = 2'b00;    end
        { 4'b1010 , 4'b0001 , 1'b1 }: begin     s = 4'b1100;    co = 2'b00;    end
        { 4'b1010 , 4'b0010 , 1'b0 }: begin     s = 4'b1100;    co = 2'b00;    end
        { 4'b1010 , 4'b0010 , 1'b1 }: begin     s = 4'b1101;    co = 2'b00;    end
        { 4'b1010 , 4'b0011 , 1'b0 }: begin     s = 4'b1101;    co = 2'b00;    end
        { 4'b1010 , 4'b0011 , 1'b1 }: begin     s = 4'b1110;    co = 2'b00;    end
        { 4'b1010 , 4'b0100 , 1'b0 }: begin     s = 4'b1110;    co = 2'b00;    end
        { 4'b1010 , 4'b0100 , 1'b1 }: begin     s = 4'b1111;    co = 2'b00;    end
        { 4'b1010 , 4'b0101 , 1'b0 }: begin     s = 4'b1111;    co = 2'b00;    end
        { 4'b1010 , 4'b0101 , 1'b1 }: begin     s = 4'b0000;    co = 2'b01;    end
        { 4'b1010 , 4'b0110 , 1'b0 }: begin     s = 4'b0000;    co = 2'b01;    end
        { 4'b1010 , 4'b0110 , 1'b1 }: begin     s = 4'b0001;    co = 2'b01;    end
        { 4'b1010 , 4'b0111 , 1'b0 }: begin     s = 4'b0001;    co = 2'b01;    end
        { 4'b1010 , 4'b0111 , 1'b1 }: begin     s = 4'b0010;    co = 2'b01;    end
        { 4'b1010 , 4'b1000 , 1'b0 }: begin     s = 4'b0010;    co = 2'b01;    end
        { 4'b1010 , 4'b1000 , 1'b1 }: begin     s = 4'b0011;    co = 2'b01;    end
        { 4'b1010 , 4'b1001 , 1'b0 }: begin     s = 4'b0011;    co = 2'b01;    end
        { 4'b1010 , 4'b1001 , 1'b1 }: begin     s = 4'b0100;    co = 2'b01;    end
        { 4'b1010 , 4'b1010 , 1'b0 }: begin     s = 4'b0100;    co = 2'b01;    end
        { 4'b1010 , 4'b1010 , 1'b1 }: begin     s = 4'b0101;    co = 2'b01;    end
        { 4'b1010 , 4'b1011 , 1'b0 }: begin     s = 4'b0101;    co = 2'b01;    end
        { 4'b1010 , 4'b1011 , 1'b1 }: begin     s = 4'b0110;    co = 2'b01;    end
        { 4'b1010 , 4'b1100 , 1'b0 }: begin     s = 4'b0110;    co = 2'b01;    end
        { 4'b1010 , 4'b1100 , 1'b1 }: begin     s = 4'b0111;    co = 2'b01;    end
        { 4'b1010 , 4'b1101 , 1'b0 }: begin     s = 4'b0111;    co = 2'b01;    end
        { 4'b1010 , 4'b1101 , 1'b1 }: begin     s = 4'b1000;    co = 2'b01;    end
        { 4'b1010 , 4'b1110 , 1'b0 }: begin     s = 4'b1000;    co = 2'b01;    end
        { 4'b1010 , 4'b1110 , 1'b1 }: begin     s = 4'b1001;    co = 2'b01;    end
        { 4'b1010 , 4'b1111 , 1'b0 }: begin     s = 4'b1001;    co = 2'b01;    end
        { 4'b1010 , 4'b1111 , 1'b1 }: begin     s = 4'b1010;    co = 2'b01;    end
        //  a=B, b=0~F, c=0~1, truth table check ( OK )
        { 4'b1011 , 4'b0000 , 1'b0 }: begin     s = 4'b1011;    co = 2'b00;    end
        { 4'b1011 , 4'b0000 , 1'b1 }: begin     s = 4'b1100;    co = 2'b00;    end
        { 4'b1011 , 4'b0001 , 1'b0 }: begin     s = 4'b1100;    co = 2'b00;    end
        { 4'b1011 , 4'b0001 , 1'b1 }: begin     s = 4'b1101;    co = 2'b00;    end
        { 4'b1011 , 4'b0010 , 1'b0 }: begin     s = 4'b1101;    co = 2'b00;    end
        { 4'b1011 , 4'b0010 , 1'b1 }: begin     s = 4'b1110;    co = 2'b00;    end
        { 4'b1011 , 4'b0011 , 1'b0 }: begin     s = 4'b1110;    co = 2'b00;    end
        { 4'b1011 , 4'b0011 , 1'b1 }: begin     s = 4'b1111;    co = 2'b00;    end
        { 4'b1011 , 4'b0100 , 1'b0 }: begin     s = 4'b1111;    co = 2'b00;    end
        { 4'b1011 , 4'b0100 , 1'b1 }: begin     s = 4'b0000;    co = 2'b01;    end
        { 4'b1011 , 4'b0101 , 1'b0 }: begin     s = 4'b0000;    co = 2'b01;    end
        { 4'b1011 , 4'b0101 , 1'b1 }: begin     s = 4'b0001;    co = 2'b01;    end
        { 4'b1011 , 4'b0110 , 1'b0 }: begin     s = 4'b0001;    co = 2'b01;    end
        { 4'b1011 , 4'b0110 , 1'b1 }: begin     s = 4'b0010;    co = 2'b01;    end
        { 4'b1011 , 4'b0111 , 1'b0 }: begin     s = 4'b0010;    co = 2'b01;    end
        { 4'b1011 , 4'b0111 , 1'b1 }: begin     s = 4'b0011;    co = 2'b01;    end
        { 4'b1011 , 4'b1000 , 1'b0 }: begin     s = 4'b0011;    co = 2'b01;    end
        { 4'b1011 , 4'b1000 , 1'b1 }: begin     s = 4'b0100;    co = 2'b01;    end
        { 4'b1011 , 4'b1001 , 1'b0 }: begin     s = 4'b0100;    co = 2'b01;    end
        { 4'b1011 , 4'b1001 , 1'b1 }: begin     s = 4'b0101;    co = 2'b01;    end
        { 4'b1011 , 4'b1010 , 1'b0 }: begin     s = 4'b0101;    co = 2'b01;    end
        { 4'b1011 , 4'b1010 , 1'b1 }: begin     s = 4'b0110;    co = 2'b01;    end
        { 4'b1011 , 4'b1011 , 1'b0 }: begin     s = 4'b0110;    co = 2'b01;    end
        { 4'b1011 , 4'b1011 , 1'b1 }: begin     s = 4'b0111;    co = 2'b01;    end
        { 4'b1011 , 4'b1100 , 1'b0 }: begin     s = 4'b0111;    co = 2'b01;    end
        { 4'b1011 , 4'b1100 , 1'b1 }: begin     s = 4'b1000;    co = 2'b01;    end
        { 4'b1011 , 4'b1101 , 1'b0 }: begin     s = 4'b1000;    co = 2'b01;    end
        { 4'b1011 , 4'b1101 , 1'b1 }: begin     s = 4'b1001;    co = 2'b01;    end
        { 4'b1011 , 4'b1110 , 1'b0 }: begin     s = 4'b1001;    co = 2'b01;    end
        { 4'b1011 , 4'b1110 , 1'b1 }: begin     s = 4'b1010;    co = 2'b01;    end
        { 4'b1011 , 4'b1111 , 1'b0 }: begin     s = 4'b1010;    co = 2'b01;    end
        { 4'b1011 , 4'b1111 , 1'b1 }: begin     s = 4'b1011;    co = 2'b01;    end
        //  a=C, b=0~F, c=0~1, truth table check ( OK )
        { 4'b1100 , 4'b0000 , 1'b0 }: begin     s = 4'b1100;    co = 2'b00;    end
        { 4'b1100 , 4'b0000 , 1'b1 }: begin     s = 4'b1101;    co = 2'b00;    end
        { 4'b1100 , 4'b0001 , 1'b0 }: begin     s = 4'b1101;    co = 2'b00;    end
        { 4'b1100 , 4'b0001 , 1'b1 }: begin     s = 4'b1110;    co = 2'b00;    end
        { 4'b1100 , 4'b0010 , 1'b0 }: begin     s = 4'b1110;    co = 2'b00;    end
        { 4'b1100 , 4'b0010 , 1'b1 }: begin     s = 4'b1111;    co = 2'b00;    end
        { 4'b1100 , 4'b0011 , 1'b0 }: begin     s = 4'b1111;    co = 2'b00;    end
        { 4'b1100 , 4'b0011 , 1'b1 }: begin     s = 4'b0000;    co = 2'b01;    end
        { 4'b1100 , 4'b0100 , 1'b0 }: begin     s = 4'b0000;    co = 2'b01;    end
        { 4'b1100 , 4'b0100 , 1'b1 }: begin     s = 4'b0001;    co = 2'b01;    end
        { 4'b1100 , 4'b0101 , 1'b0 }: begin     s = 4'b0001;    co = 2'b01;    end
        { 4'b1100 , 4'b0101 , 1'b1 }: begin     s = 4'b0010;    co = 2'b01;    end
        { 4'b1100 , 4'b0110 , 1'b0 }: begin     s = 4'b0010;    co = 2'b01;    end
        { 4'b1100 , 4'b0110 , 1'b1 }: begin     s = 4'b0011;    co = 2'b01;    end
        { 4'b1100 , 4'b0111 , 1'b0 }: begin     s = 4'b0011;    co = 2'b01;    end
        { 4'b1100 , 4'b0111 , 1'b1 }: begin     s = 4'b0100;    co = 2'b01;    end
        { 4'b1100 , 4'b1000 , 1'b0 }: begin     s = 4'b0100;    co = 2'b01;    end
        { 4'b1100 , 4'b1000 , 1'b1 }: begin     s = 4'b0101;    co = 2'b01;    end
        { 4'b1100 , 4'b1001 , 1'b0 }: begin     s = 4'b0101;    co = 2'b01;    end
        { 4'b1100 , 4'b1001 , 1'b1 }: begin     s = 4'b0110;    co = 2'b01;    end
        { 4'b1100 , 4'b1010 , 1'b0 }: begin     s = 4'b0110;    co = 2'b01;    end
        { 4'b1100 , 4'b1010 , 1'b1 }: begin     s = 4'b0111;    co = 2'b01;    end
        { 4'b1100 , 4'b1011 , 1'b0 }: begin     s = 4'b0111;    co = 2'b01;    end
        { 4'b1100 , 4'b1011 , 1'b1 }: begin     s = 4'b1000;    co = 2'b01;    end
        { 4'b1100 , 4'b1100 , 1'b0 }: begin     s = 4'b1000;    co = 2'b01;    end
        { 4'b1100 , 4'b1100 , 1'b1 }: begin     s = 4'b1001;    co = 2'b01;    end
        { 4'b1100 , 4'b1101 , 1'b0 }: begin     s = 4'b1001;    co = 2'b01;    end
        { 4'b1100 , 4'b1101 , 1'b1 }: begin     s = 4'b1010;    co = 2'b01;    end
        { 4'b1100 , 4'b1110 , 1'b0 }: begin     s = 4'b1010;    co = 2'b01;    end
        { 4'b1100 , 4'b1110 , 1'b1 }: begin     s = 4'b1011;    co = 2'b01;    end
        { 4'b1100 , 4'b1111 , 1'b0 }: begin     s = 4'b1011;    co = 2'b01;    end
        { 4'b1100 , 4'b1111 , 1'b1 }: begin     s = 4'b1100;    co = 2'b01;    end
        //  a=D, b=0~F, c=0~1, truth table check ( OK )
        { 4'b1101 , 4'b0000 , 1'b0 }: begin     s = 4'b1101;    co = 2'b00;    end
        { 4'b1101 , 4'b0000 , 1'b1 }: begin     s = 4'b1110;    co = 2'b00;    end
        { 4'b1101 , 4'b0001 , 1'b0 }: begin     s = 4'b1110;    co = 2'b00;    end
        { 4'b1101 , 4'b0001 , 1'b1 }: begin     s = 4'b1111;    co = 2'b00;    end
        { 4'b1101 , 4'b0010 , 1'b0 }: begin     s = 4'b1111;    co = 2'b00;    end
        { 4'b1101 , 4'b0010 , 1'b1 }: begin     s = 4'b0000;    co = 2'b01;    end
        { 4'b1101 , 4'b0011 , 1'b0 }: begin     s = 4'b0000;    co = 2'b01;    end
        { 4'b1101 , 4'b0011 , 1'b1 }: begin     s = 4'b0001;    co = 2'b01;    end
        { 4'b1101 , 4'b0100 , 1'b0 }: begin     s = 4'b0001;    co = 2'b01;    end
        { 4'b1101 , 4'b0100 , 1'b1 }: begin     s = 4'b0010;    co = 2'b01;    end
        { 4'b1101 , 4'b0101 , 1'b0 }: begin     s = 4'b0010;    co = 2'b01;    end
        { 4'b1101 , 4'b0101 , 1'b1 }: begin     s = 4'b0011;    co = 2'b01;    end
        { 4'b1101 , 4'b0110 , 1'b0 }: begin     s = 4'b0011;    co = 2'b01;    end
        { 4'b1101 , 4'b0110 , 1'b1 }: begin     s = 4'b0100;    co = 2'b01;    end
        { 4'b1101 , 4'b0111 , 1'b0 }: begin     s = 4'b0100;    co = 2'b01;    end
        { 4'b1101 , 4'b0111 , 1'b1 }: begin     s = 4'b0101;    co = 2'b01;    end
        { 4'b1101 , 4'b1000 , 1'b0 }: begin     s = 4'b0101;    co = 2'b01;    end
        { 4'b1101 , 4'b1000 , 1'b1 }: begin     s = 4'b0110;    co = 2'b01;    end
        { 4'b1101 , 4'b1001 , 1'b0 }: begin     s = 4'b0110;    co = 2'b01;    end
        { 4'b1101 , 4'b1001 , 1'b1 }: begin     s = 4'b0111;    co = 2'b01;    end
        { 4'b1101 , 4'b1010 , 1'b0 }: begin     s = 4'b0111;    co = 2'b01;    end
        { 4'b1101 , 4'b1010 , 1'b1 }: begin     s = 4'b1000;    co = 2'b01;    end
        { 4'b1101 , 4'b1011 , 1'b0 }: begin     s = 4'b1000;    co = 2'b01;    end
        { 4'b1101 , 4'b1011 , 1'b1 }: begin     s = 4'b1001;    co = 2'b01;    end
        { 4'b1101 , 4'b1100 , 1'b0 }: begin     s = 4'b1001;    co = 2'b01;    end
        { 4'b1101 , 4'b1100 , 1'b1 }: begin     s = 4'b1010;    co = 2'b01;    end
        { 4'b1101 , 4'b1101 , 1'b0 }: begin     s = 4'b1010;    co = 2'b01;    end
        { 4'b1101 , 4'b1101 , 1'b1 }: begin     s = 4'b1011;    co = 2'b01;    end
        { 4'b1101 , 4'b1110 , 1'b0 }: begin     s = 4'b1011;    co = 2'b01;    end
        { 4'b1101 , 4'b1110 , 1'b1 }: begin     s = 4'b1100;    co = 2'b01;    end
        { 4'b1101 , 4'b1111 , 1'b0 }: begin     s = 4'b1100;    co = 2'b01;    end
        { 4'b1101 , 4'b1111 , 1'b1 }: begin     s = 4'b1101;    co = 2'b01;    end
        //  a=E, b=0~F, c=0~1, truth table check ( OK )
        { 4'b1110 , 4'b0000 , 1'b0 }: begin     s = 4'b1110;    co = 2'b00;    end
        { 4'b1110 , 4'b0000 , 1'b1 }: begin     s = 4'b1111;    co = 2'b00;    end
        { 4'b1110 , 4'b0001 , 1'b0 }: begin     s = 4'b1111;    co = 2'b00;    end
        { 4'b1110 , 4'b0001 , 1'b1 }: begin     s = 4'b0000;    co = 2'b01;    end
        { 4'b1110 , 4'b0010 , 1'b0 }: begin     s = 4'b0000;    co = 2'b01;    end
        { 4'b1110 , 4'b0010 , 1'b1 }: begin     s = 4'b0001;    co = 2'b01;    end
        { 4'b1110 , 4'b0011 , 1'b0 }: begin     s = 4'b0001;    co = 2'b01;    end
        { 4'b1110 , 4'b0011 , 1'b1 }: begin     s = 4'b0010;    co = 2'b01;    end
        { 4'b1110 , 4'b0100 , 1'b0 }: begin     s = 4'b0010;    co = 2'b01;    end
        { 4'b1110 , 4'b0100 , 1'b1 }: begin     s = 4'b0011;    co = 2'b01;    end
        { 4'b1110 , 4'b0101 , 1'b0 }: begin     s = 4'b0011;    co = 2'b01;    end
        { 4'b1110 , 4'b0101 , 1'b1 }: begin     s = 4'b0100;    co = 2'b01;    end
        { 4'b1110 , 4'b0110 , 1'b0 }: begin     s = 4'b0100;    co = 2'b01;    end
        { 4'b1110 , 4'b0110 , 1'b1 }: begin     s = 4'b0101;    co = 2'b01;    end
        { 4'b1110 , 4'b0111 , 1'b0 }: begin     s = 4'b0101;    co = 2'b01;    end
        { 4'b1110 , 4'b0111 , 1'b1 }: begin     s = 4'b0110;    co = 2'b01;    end
        { 4'b1110 , 4'b1000 , 1'b0 }: begin     s = 4'b0110;    co = 2'b01;    end
        { 4'b1110 , 4'b1000 , 1'b1 }: begin     s = 4'b0111;    co = 2'b01;    end
        { 4'b1110 , 4'b1001 , 1'b0 }: begin     s = 4'b0111;    co = 2'b01;    end
        { 4'b1110 , 4'b1001 , 1'b1 }: begin     s = 4'b1000;    co = 2'b01;    end
        { 4'b1110 , 4'b1010 , 1'b0 }: begin     s = 4'b1000;    co = 2'b01;    end
        { 4'b1110 , 4'b1010 , 1'b1 }: begin     s = 4'b1001;    co = 2'b01;    end
        { 4'b1110 , 4'b1011 , 1'b0 }: begin     s = 4'b1001;    co = 2'b01;    end
        { 4'b1110 , 4'b1011 , 1'b1 }: begin     s = 4'b1010;    co = 2'b01;    end
        { 4'b1110 , 4'b1100 , 1'b0 }: begin     s = 4'b1010;    co = 2'b01;    end
        { 4'b1110 , 4'b1100 , 1'b1 }: begin     s = 4'b1011;    co = 2'b01;    end
        { 4'b1110 , 4'b1101 , 1'b0 }: begin     s = 4'b1011;    co = 2'b01;    end
        { 4'b1110 , 4'b1101 , 1'b1 }: begin     s = 4'b1100;    co = 2'b01;    end
        { 4'b1110 , 4'b1110 , 1'b0 }: begin     s = 4'b1100;    co = 2'b01;    end
        { 4'b1110 , 4'b1110 , 1'b1 }: begin     s = 4'b1101;    co = 2'b01;    end
        { 4'b1110 , 4'b1111 , 1'b0 }: begin     s = 4'b1101;    co = 2'b01;    end
        { 4'b1110 , 4'b1111 , 1'b1 }: begin     s = 4'b1110;    co = 2'b10;    end
        //  a=F, b=0~F, c=0~1, truth table check ( OK )
        { 4'b1111 , 4'b0000 , 1'b0 }: begin     s = 4'b1111;    co = 2'b00;    end
        { 4'b1111 , 4'b0000 , 1'b1 }: begin     s = 4'b0000;    co = 2'b01;    end
        { 4'b1111 , 4'b0001 , 1'b0 }: begin     s = 4'b0000;    co = 2'b01;    end
        { 4'b1111 , 4'b0001 , 1'b1 }: begin     s = 4'b0001;    co = 2'b01;    end
        { 4'b1111 , 4'b0010 , 1'b0 }: begin     s = 4'b0001;    co = 2'b01;    end
        { 4'b1111 , 4'b0010 , 1'b1 }: begin     s = 4'b0010;    co = 2'b01;    end
        { 4'b1111 , 4'b0011 , 1'b0 }: begin     s = 4'b0010;    co = 2'b01;    end
        { 4'b1111 , 4'b0011 , 1'b1 }: begin     s = 4'b0011;    co = 2'b01;    end
        { 4'b1111 , 4'b0100 , 1'b0 }: begin     s = 4'b0011;    co = 2'b01;    end
        { 4'b1111 , 4'b0100 , 1'b1 }: begin     s = 4'b0100;    co = 2'b01;    end
        { 4'b1111 , 4'b0101 , 1'b0 }: begin     s = 4'b0100;    co = 2'b01;    end
        { 4'b1111 , 4'b0101 , 1'b1 }: begin     s = 4'b0101;    co = 2'b01;    end
        { 4'b1111 , 4'b0110 , 1'b0 }: begin     s = 4'b0101;    co = 2'b01;    end
        { 4'b1111 , 4'b0110 , 1'b1 }: begin     s = 4'b0110;    co = 2'b01;    end
        { 4'b1111 , 4'b0111 , 1'b0 }: begin     s = 4'b0110;    co = 2'b01;    end
        { 4'b1111 , 4'b0111 , 1'b1 }: begin     s = 4'b0111;    co = 2'b01;    end
        { 4'b1111 , 4'b1000 , 1'b0 }: begin     s = 4'b0111;    co = 2'b01;    end
        { 4'b1111 , 4'b1000 , 1'b1 }: begin     s = 4'b1000;    co = 2'b01;    end
        { 4'b1111 , 4'b1001 , 1'b0 }: begin     s = 4'b1000;    co = 2'b01;    end
        { 4'b1111 , 4'b1001 , 1'b1 }: begin     s = 4'b1001;    co = 2'b01;    end
        { 4'b1111 , 4'b1010 , 1'b0 }: begin     s = 4'b1001;    co = 2'b01;    end
        { 4'b1111 , 4'b1010 , 1'b1 }: begin     s = 4'b1010;    co = 2'b01;    end
        { 4'b1111 , 4'b1011 , 1'b0 }: begin     s = 4'b1010;    co = 2'b01;    end
        { 4'b1111 , 4'b1011 , 1'b1 }: begin     s = 4'b1011;    co = 2'b01;    end
        { 4'b1111 , 4'b1100 , 1'b0 }: begin     s = 4'b1011;    co = 2'b01;    end
        { 4'b1111 , 4'b1100 , 1'b1 }: begin     s = 4'b1100;    co = 2'b01;    end
        { 4'b1111 , 4'b1101 , 1'b0 }: begin     s = 4'b1100;    co = 2'b01;    end
        { 4'b1111 , 4'b1101 , 1'b1 }: begin     s = 4'b1101;    co = 2'b01;    end
        { 4'b1111 , 4'b1110 , 1'b0 }: begin     s = 4'b1101;    co = 2'b01;    end
        { 4'b1111 , 4'b1110 , 1'b1 }: begin     s = 4'b1110;    co = 2'b10;    end
        { 4'b1111 , 4'b1111 , 1'b0 }: begin     s = 4'b1110;    co = 2'b10;    end
        { 4'b1111 , 4'b1111 , 1'b1 }: begin     s = 4'b1111;    co = 2'b10;    end
        endcase
    end
endmodule
