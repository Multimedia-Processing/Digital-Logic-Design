module or_gate (a,b,c);

input a,b;
output c;
or(a,b,c);
    
endmodule