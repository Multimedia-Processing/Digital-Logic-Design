
`timescale 1ns/1ps

module T;
    reg [3:0] D0 = 4'b0101;
    reg [3:0] D1 = 4'b1111;
    reg [3:0] D2 = 4'b1111;
    reg [3:0] D3 = 4'b0101;
    reg [1:0] S = 2'b00;
    wire [3:0] Y;


    mux4_1 UUT (
        .D0(D0),
        .D1(D1),
        .D2(D2),
        .D3(D3),
        .S(S),
        .Y(Y));

    initial
    begin
      #2000 // Final time:  2000 ns
        $stop;
    end

    initial begin
        // -------------  Current Time:  100ns
        #100;
        D0 = 4'b1100;
        D1 = 4'b1010;
        D2 = 4'b0010;
        D3 = 4'b1001;
        // -------------------------------------
        // -------------  Current Time:  200ns
        #100;
        D0 = 4'b1001;
        D1 = 4'b0000;
        D2 = 4'b1010;
        D3 = 4'b1000;
        // -------------------------------------
        // -------------  Current Time:  300ns
        #100;
        D0 = 4'b0001;
        D1 = 4'b1001;
        D2 = 4'b1111;
        D3 = 4'b0111;
        // -------------------------------------
        // -------------  Current Time:  400ns
        #100;
        D0 = 4'b1110;
        D1 = 4'b0100;
        D2 = 4'b0110;
        D3 = 4'b1111;
        // -------------------------------------
        // -------------  Current Time:  500ns
        #100;
        D0 = 4'b0111;
        D1 = 4'b0101;
        D2 = 4'b1100;
        D3 = 4'b0110;
        S = 2'b01;
        // -------------------------------------
        // -------------  Current Time:  600ns
        #100;
        D0 = 4'b1000;
        D1 = 4'b1001;
        D2 = 4'b0001;
        D3 = 4'b0011;
        // -------------------------------------
        // -------------  Current Time:  700ns
        #100;
        D0 = 4'b1010;
        D1 = 4'b0000;
        D2 = 4'b0000;
        D3 = 4'b1011;
        // -------------------------------------
        // -------------  Current Time:  800ns
        #100;
        D0 = 4'b0011;
        D1 = 4'b0011;
        D2 = 4'b1100;
        D3 = 4'b0100;
        // -------------------------------------
        // -------------  Current Time:  900ns
        #100;
        D0 = 4'b0110;
        D1 = 4'b1111;
        D2 = 4'b0101;
        D3 = 4'b1101;
        // -------------------------------------
        // -------------  Current Time:  1000ns
        #100;
        D0 = 4'b1100;
        D1 = 4'b0110;
        D2 = 4'b1100;
        D3 = 4'b1001;
        S = 2'b10;
        // -------------------------------------
        // -------------  Current Time:  1100ns
        #100;
        D0 = 4'b0001;
        D1 = 4'b1011;
        D2 = 4'b1010;
        D3 = 4'b0000;
        // -------------------------------------
        // -------------  Current Time:  1200ns
        #100;
        D0 = 4'b1000;
        D1 = 4'b1100;
        D2 = 4'b0011;
        D3 = 4'b1001;
        // -------------------------------------
        // -------------  Current Time:  1300ns
        #100;
        D0 = 4'b1001;
        D1 = 4'b0000;
        D2 = 4'b1110;
        D3 = 4'b1101;
        // -------------------------------------
        // -------------  Current Time:  1400ns
        #100;
        D0 = 4'b0101;
        D1 = 4'b1101;
        D2 = 4'b0110;
        D3 = 4'b0110;
        // -------------------------------------
        // -------------  Current Time:  1500ns
        #100;
        D0 = 4'b1100;
        D1 = 4'b0101;
        D2 = 4'b0111;
        D3 = 4'b1011;
        S = 2'b11;
        // -------------------------------------
        // -------------  Current Time:  1600ns
        #100;
        D0 = 4'b0010;
        D1 = 4'b0000;
        D2 = 4'b1010;
        D3 = 4'b0010;
        // -------------------------------------
        // -------------  Current Time:  1700ns
        #100;
        D0 = 4'b0011;
        D1 = 4'b1001;
        D2 = 4'b0000;
        D3 = 4'b0001;
        // -------------------------------------
        // -------------  Current Time:  1800ns
        #100;
        D0 = 4'b1010;
        D1 = 4'b0001;
        D2 = 4'b0101;
        D3 = 4'b1111;
        // -------------------------------------
        // -------------  Current Time:  1900ns
        #100;
        D0 = 4'b0110;
        D1 = 4'b1110;
        D2 = 4'b1100;
        D3 = 4'b0110;
    end

endmodule

