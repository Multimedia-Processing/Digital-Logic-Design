module and_date (a, b, c);
input a, b;
output c;

assign c = a & b;

endmodule // and_date
