module snake ();

endmodule // snake
