module nor_gate(a,b,nor_output);

input a,b;
output nor_output;
nor(nor_output,a,b);

endmodule
