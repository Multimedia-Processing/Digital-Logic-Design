////////////////////////////////////////////////////////////////////////////////

`timescale 1ns/1ps

module T;
    reg [2:0] S = 3'b000;
    reg [3:0] A = 4'b0000;
    reg [3:0] B = 4'b1111;
    wire [4:0] Alu1;
    wire [4:0] Alu2;


    alu4 UUT (
        .S(S),
        .A(A),
        .B(B),
        .Alu1(Alu1),
        .Alu2(Alu2));

    initial
    begin
      #4000 // Final time:  4000 ns
        $stop;
    end

    initial begin
        // -------------  Current Time:  100ns
        #100;
        A = 4'b1000;
        B = 4'b0010;
        // -------------------------------------
        // -------------  Current Time:  200ns
        #100;
        A = 4'b1001;
        B = 4'b0011;
        // -------------------------------------
        // -------------  Current Time:  300ns
        #100;
        A = 4'b0001;
        B = 4'b1110;
        // -------------------------------------
        // -------------  Current Time:  400ns
        #100;
        A = 4'b1110;
        B = 4'b0110;
        // -------------------------------------
        // -------------  Current Time:  500ns
        #100;
        A = 4'b0111;
        B = 4'b0111;
        S = 3'b001;
        // -------------------------------------
        // -------------  Current Time:  600ns
        #100;
        B = 4'b1010;
        // -------------------------------------
        // -------------  Current Time:  700ns
        #100;
        A = 4'b1010;
        B = 4'b0000;
        // -------------------------------------
        // -------------  Current Time:  800ns
        #100;
        A = 4'b0011;
        B = 4'b0101;
        // -------------------------------------
        // -------------  Current Time:  900ns
        #100;
        A = 4'b0110;
        B = 4'b1100;
        // -------------------------------------
        // -------------  Current Time:  1000ns
        #100;
        A = 4'b1100;
        B = 4'b0101;
        S = 3'b010;
        // -------------------------------------
        // -------------  Current Time:  1100ns
        #100;
        A = 4'b0001;
        B = 4'b1001;
        // -------------------------------------
        // -------------  Current Time:  1200ns
        #100;
        A = 4'b1000;
        B = 4'b1000;
        // -------------------------------------
        // -------------  Current Time:  1300ns
        #100;
        B = 4'b0111;
        // -------------------------------------
        // -------------  Current Time:  1400ns
        #100;
        A = 4'b0101;
        B = 4'b1111;
        // -------------------------------------
        // -------------  Current Time:  1500ns
        #100;
        A = 4'b1100;
        B = 4'b0110;
        S = 3'b100;
        // -------------------------------------
        // -------------  Current Time:  1600ns
        #100;
        A = 4'b0010;
        B = 4'b0011;
        // -------------------------------------
        // -------------  Current Time:  1700ns
        #100;
        A = 4'b0011;
        B = 4'b1011;
        // -------------------------------------
        // -------------  Current Time:  1800ns
        #100;
        A = 4'b1010;
        B = 4'b0100;
        // -------------------------------------
        // -------------  Current Time:  1900ns
        #100;
        A = 4'b0110;
        B = 4'b1101;
        // -------------------------------------
        // -------------  Current Time:  2000ns
        #100;
        A = 4'b1111;
        B = 4'b1001;
        S = 3'b011;
        // -------------------------------------
        // -------------  Current Time:  2100ns
        #100;
        A = 4'b1010;
        B = 4'b0000;
        // -------------------------------------
        // -------------  Current Time:  2200ns
        #100;
        A = 4'b0000;
        B = 4'b1001;
        S = 3'b101;
        // -------------------------------------
        // -------------  Current Time:  2300ns
        #100;
        A = 4'b1001;
        B = 4'b1101;
        // -------------------------------------
        // -------------  Current Time:  2400ns
        #100;
        A = 4'b0100;
        B = 4'b0110;
        S = 3'b110;
        // -------------------------------------
        // -------------  Current Time:  2500ns
        #100;
        A = 4'b0101;
        B = 4'b1011;
        // -------------------------------------
        // -------------  Current Time:  2600ns
        #100;
        A = 4'b1001;
        B = 4'b0010;
        S = 3'b111;
        // -------------------------------------
        // -------------  Current Time:  2700ns
        #100;
        A = 4'b0000;
        // -------------------------------------
        // -------------  Current Time:  2800ns
        #100;
        A = 4'b0011;
        B = 4'b1111;
        // -------------------------------------
        // -------------  Current Time:  2900ns
        #100;
        A = 4'b1111;
        B = 4'b0110;
        // -------------------------------------
        // -------------  Current Time:  3000ns
        #100;
        A = 4'b0110;
        B = 4'b1000;
        // -------------------------------------
        // -------------  Current Time:  3100ns
        #100;
        A = 4'b1011;
        B = 4'b1001;
        // -------------------------------------
        // -------------  Current Time:  3200ns
        #100;
        B = 4'b0000;
        // -------------------------------------
        // -------------  Current Time:  3300ns
        #100;
        A = 4'b0000;
        B = 4'b1100;
        // -------------------------------------
        // -------------  Current Time:  3400ns
        #100;
        A = 4'b1101;
        B = 4'b0101;
        // -------------------------------------
        // -------------  Current Time:  3500ns
        #100;
        A = 4'b0101;
        B = 4'b0000;
        // -------------------------------------
        // -------------  Current Time:  3600ns
        #100;
        A = 4'b0000;
        B = 4'b1010;
        // -------------------------------------
        // -------------  Current Time:  3700ns
        #100;
        A = 4'b1001;
        B = 4'b0011;
        // -------------------------------------
        // -------------  Current Time:  3800ns
        #100;
        A = 4'b0001;
        B = 4'b1110;
        // -------------------------------------
        // -------------  Current Time:  3900ns
        #100;
        A = 4'b1110;
        // -------------------------------------
        // -------------  Current Time:  4000ns
        #100;
        A = 4'b1111;
        B = 4'b0011;
    end

endmodule

