module and_gate(a,b,o);
input a,b;
output o;

and (o,a,b);


endmodule