module not_gate (a, b, c, d);

input a, b;
output c, d;
not(c, a);
not(d, b);
    
endmodule