module arithmetic_logic_shift_unit(
    operation_select,
    operation,
    function_output
);
