
`timescale 1ns/1ps

module T;
    reg [3:0] A = 4'b0000;
    reg [3:0] B = 4'b0000;
    reg Ci = 1'b0;
    wire Co;
    wire [3:0] S;
    wire [3:0] X;
    wire [3:0] Y;
    wire [3:0] Z;


    op UUT (
        .A(A),
        .B(B),
        .Ci(Ci),
        .Co(Co),
        .S(S),
        .X(X),
        .Y(Y),
        .Z(Z));

    initial
    begin
      #1000 // Final time:  1000 ns
        $stop;
    end

    initial begin
        // -------------  Current Time:  100ns
        #100;
        Ci = 1'b1;
        A = 4'b1100;
        B = 4'b1010;
        // -------------------------------------
        // -------------  Current Time:  200ns
        #100;
        Ci = 1'b0;
        A = 4'b1001;
        B = 4'b0000;
        // -------------------------------------
        // -------------  Current Time:  300ns
        #100;
        Ci = 1'b1;
        A = 4'b0001;
        B = 4'b1001;
        // -------------------------------------
        // -------------  Current Time:  400ns
        #100;
        Ci = 1'b0;
        A = 4'b1110;
        B = 4'b0100;
        // -------------------------------------
        // -------------  Current Time:  500ns
        #100;
        Ci = 1'b1;
        A = 4'b0111;
        B = 4'b0101;
        // -------------------------------------
        // -------------  Current Time:  600ns
        #100;
        Ci = 1'b0;
        A = 4'b1000;
        B = 4'b1001;
        // -------------------------------------
        // -------------  Current Time:  700ns
        #100;
        Ci = 1'b1;
        A = 4'b1010;
        B = 4'b0000;
        // -------------------------------------
        // -------------  Current Time:  800ns
        #100;
        Ci = 1'b0;
        A = 4'b0011;
        B = 4'b0011;
        // -------------------------------------
        // -------------  Current Time:  900ns
        #100;
        Ci = 1'b1;
        A = 4'b1111;
        B = 4'b1111;
        // -------------------------------------
        // -------------  Current Time:  1000ns
        #100;
        A = 4'b1101;
        B = 4'b0110;
    end

endmodule

