////////////////////////////////////////////////////////////////////////////////

`timescale 1ns/1ps

module T;
    reg Clk = 1'b0;
    reg [3:0] D = 4'b0101;
    wire [3:0] Q_l;
    wire [3:0] Q_ff;


    d_latch_ff UUT (
        .Clk(Clk),
        .D(D),
        .Q_l(Q_l),
        .Q_ff(Q_ff));

    initial
    begin
      #2000 // Final time:  2000 ns
        $stop;
    end

    initial begin
        // -------------  Current Time:  100ns
        #100;
        Clk = 1'b1;
        D = 4'b1100;
        // -------------------------------------
        // -------------  Current Time:  200ns
        #100;
        D = 4'b1001;
        // -------------------------------------
        // -------------  Current Time:  300ns
        #100;
        Clk = 1'b0;
        D = 4'b0001;
        // -------------------------------------
        // -------------  Current Time:  400ns
        #100;
        D = 4'b1110;
        // -------------------------------------
        // -------------  Current Time:  500ns
        #100;
        Clk = 1'b1;
        D = 4'b0111;
        // -------------------------------------
        // -------------  Current Time:  600ns
        #100;
        D = 4'b1001;
        // -------------------------------------
        // -------------  Current Time:  700ns
        #100;
        Clk = 1'b0;
        D = 4'b1010;
        // -------------------------------------
        // -------------  Current Time:  800ns
        #100;
        D = 4'b0011;
        // -------------------------------------
        // -------------  Current Time:  900ns
        #100;
        Clk = 1'b1;
        D = 4'b0110;
        // -------------------------------------
        // -------------  Current Time:  1000ns
        #100;
        D = 4'b1100;
        // -------------------------------------
        // -------------  Current Time:  1100ns
        #100;
        Clk = 1'b0;
        D = 4'b0001;
        // -------------------------------------
        // -------------  Current Time:  1200ns
        #100;
        D = 4'b1000;
        // -------------------------------------
        // -------------  Current Time:  1300ns
        #100;
        Clk = 1'b1;
        D = 4'b0000;
        // -------------------------------------
        // -------------  Current Time:  1400ns
        #100;
        D = 4'b0101;
        // -------------------------------------
        // -------------  Current Time:  1500ns
        #100;
        Clk = 1'b0;
        D = 4'b1100;
        // -------------------------------------
        // -------------  Current Time:  1600ns
        #100;
        D = 4'b0010;
        // -------------------------------------
        // -------------  Current Time:  1700ns
        #100;
        Clk = 1'b1;
        D = 4'b0011;
        // -------------------------------------
        // -------------  Current Time:  1800ns
        #100;
        D = 4'b1010;
        // -------------------------------------
        // -------------  Current Time:  1900ns
        #100;
        Clk = 1'b0;
        D = 4'b0110;
    end

endmodule

