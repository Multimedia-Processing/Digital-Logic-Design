module NOT_GATE (c, a);

input a;
output c;

    not(c, a);

endmodule