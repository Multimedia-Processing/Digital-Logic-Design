
`timescale 1ns/1ps

module T;
    reg [7:0] D = 8'b00000001;
    wire [2:0] Q1;
    wire [2:0] Q2;

    enc83_priority UUT (
        .D(D),
        .Q1(Q1),
        .Q2(Q2));

    initial
    begin
      #2000 // Final time:  2000 ns
        $stop;
    end

    initial begin
        // -------------  Current Time:  100ns
        #100;
        D = 8'b00000010;
        // -------------------------------------
        // -------------  Current Time:  200ns
        #100;
        D = 8'b00000100;
        // -------------------------------------
        // -------------  Current Time:  300ns
        #100;
        D = 8'b00001000;
        // -------------------------------------
        // -------------  Current Time:  400ns
        #100;
        D = 8'b00010000;
        // -------------------------------------
        // -------------  Current Time:  500ns
        #100;
        D = 8'b00100000;
        // -------------------------------------
        // -------------  Current Time:  600ns
        #100;
        D = 8'b01000000;
        // -------------------------------------
        // -------------  Current Time:  700ns
        #100;
        D = 8'b10000000;
        // -------------------------------------
        // -------------  Current Time:  800ns
        #100;
        D = 8'b00110011;
        // -------------------------------------
        // -------------  Current Time:  900ns
        #100;
        D = 8'b11110110;
        // -------------------------------------
        // -------------  Current Time:  1000ns
        #100;
        D = 8'b10100100;
        // -------------------------------------
        // -------------  Current Time:  1100ns
        #100;
        D = 8'b11001000;
        // -------------------------------------
        // -------------  Current Time:  1200ns
        #100;
        D = 8'b10011000;
        // -------------------------------------
        // -------------  Current Time:  1300ns
        #100;
        D = 8'b00110000;
        // -------------------------------------
        // -------------  Current Time:  1400ns
        #100;
        D = 8'b11100000;
        // -------------------------------------
        // -------------  Current Time:  1500ns
        #100;
        D = 8'b01000000;
        // -------------------------------------
        // -------------  Current Time:  1600ns
        #100;
        D = 8'b10000000;
        // -------------------------------------
        // -------------  Current Time:  1700ns
        #100;
        D = 8'b11101100;
        // -------------------------------------
        // -------------  Current Time:  1800ns
        #100;
        D = 8'b01101011;
        // -------------------------------------
        // -------------  Current Time:  1900ns
        #100;
        D = 8'b01111010;
    end

endmodule

