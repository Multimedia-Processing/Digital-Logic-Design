module xnor_gate (a, b, c);

  input a, b ;
  output c ;

  xnor (c, a, b);

endmodule // xnor_gate
