
`timescale 1ns/1ps

module T;
    reg [7:0] D = 8'b00000001;
    wire [2:0] Q;


    enc83_case UUT (
        .D(D),
        .Q(Q));

    initial
    begin
      #1000 // Final time:  1000 ns
        $stop;
    end

    initial begin
        // -------------  Current Time:  100ns
        #100;
        D = 8'b00000010;
        // -------------------------------------
        // -------------  Current Time:  200ns
        #100;
        D = 8'b00000100;
        // -------------------------------------
        // -------------  Current Time:  300ns
        #100;
        D = 8'b00001000;
        // -------------------------------------
        // -------------  Current Time:  400ns
        #100;
        D = 8'b00010000;
        // -------------------------------------
        // -------------  Current Time:  500ns
        #100;
        D = 8'b00100000;
        // -------------------------------------
        // -------------  Current Time:  600ns
        #100;
        D = 8'b01000000;
        // -------------------------------------
        // -------------  Current Time:  700ns
        #100;
        D = 8'b10000000;
        // -------------------------------------
        // -------------  Current Time:  800ns
        #100;
        D = 8'b00000000;
    end

endmodule

