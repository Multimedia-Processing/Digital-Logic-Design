module not_gate (a, c);

  input a ;
  output c ;

  not (c, a);

endmodule // not_gate
