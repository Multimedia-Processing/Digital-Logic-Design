module nor_gate (A,B,C);
    input A,B;
    output C;
    
    nor(C,A,B);
    
endmodule