module not_gate(a,b,not_output);

input a,b;
output not_output;
nor(not_output,a,b);

endmodule
