library verilog;
use verilog.vl_types.all;
entity BCD_adder_1D_G_vlg_vec_tst is
end BCD_adder_1D_G_vlg_vec_tst;
