module XNOR_GATE (c, a, b);

input a, b;
output c;

    xnor(c, a, b);

endmodule