module adder_4_assign (a, b, s);
input signed [7:0] a, b;
output signed [8:0] s;

assign s1 = a + b;

endmodule // adder_4_assign
