module BUF_GATE_B (c, b);

input b;
output c;

    and(c, b);

endmodule