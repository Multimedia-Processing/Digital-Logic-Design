module sub_5_assign (a, b, s);
input [4:0] a, b;
output [4:0] s;

assign s = a - b;

endmodule // sub_5_assign
