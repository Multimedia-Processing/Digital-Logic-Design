module OR_GATE (c, a, b);

input a, b;
output c;

    or(c, a, b);

endmodule