module nand_gate(a,b,nand_output);

input a,b;
output nand_output;
nand(nand_output,a,b);

endmodule
