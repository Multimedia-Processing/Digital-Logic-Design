module and_gate (a,b,c);
    //輸入輸出
    input a, b;
    output c;

    and(c, a, b);

endmodule