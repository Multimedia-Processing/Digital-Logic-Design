module NOT_GATE_B (c, b);

input b;
output c;

    not(c, b);

endmodule