
`timescale 1ns/1ps

module T;
    wire [3:0] A1;
    wire [3:0] A2;
    wire [3:0] B1;
    wire [3:0] B2;
    wire [3:0] C1;
    wire [3:0] C2;
    wire [3:0] D1;
    wire [3:0] D2;
    reg [1:0] S = 2'b00;
    reg [3:0] Y = 4'b0101;


    demux UUT (
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .B2(B2),
        .C1(C1),
        .C2(C2),
        .D1(D1),
        .D2(D2),
        .S(S),
        .Y(Y));

    initial
    begin
      #2000 // Final time:  2000 ns
        $stop;
    end

    initial begin
        // -------------  Current Time:  100ns
        #100;
        Y = 4'b1100;
        // -------------------------------------
        // -------------  Current Time:  200ns
        #100;
        Y = 4'b1001;
        // -------------------------------------
        // -------------  Current Time:  300ns
        #100;
        Y = 4'b0001;
        // -------------------------------------
        // -------------  Current Time:  400ns
        #100;
        Y = 4'b1110;
        // -------------------------------------
        // -------------  Current Time:  500ns
        #100;
        S = 2'b01;
        Y = 4'b0111;
        // -------------------------------------
        // -------------  Current Time:  600ns
        #100;
        Y = 4'b0101;
        // -------------------------------------
        // -------------  Current Time:  700ns
        #100;
        Y = 4'b1010;
        // -------------------------------------
        // -------------  Current Time:  800ns
        #100;
        Y = 4'b0011;
        // -------------------------------------
        // -------------  Current Time:  900ns
        #100;
        Y = 4'b0110;
        // -------------------------------------
        // -------------  Current Time:  1000ns
        #100;
        S = 2'b10;
        Y = 4'b1100;
        // -------------------------------------
        // -------------  Current Time:  1100ns
        #100;
        Y = 4'b0001;
        // -------------------------------------
        // -------------  Current Time:  1200ns
        #100;
        Y = 4'b1000;
        // -------------------------------------
        // -------------  Current Time:  1300ns
        #100;
        Y = 4'b0000;
        // -------------------------------------
        // -------------  Current Time:  1400ns
        #100;
        Y = 4'b0101;
        // -------------------------------------
        // -------------  Current Time:  1500ns
        #100;
        S = 2'b11;
        Y = 4'b1100;
        // -------------------------------------
        // -------------  Current Time:  1600ns
        #100;
        Y = 4'b0010;
        // -------------------------------------
        // -------------  Current Time:  1700ns
        #100;
        Y = 4'b0011;
        // -------------------------------------
        // -------------  Current Time:  1800ns
        #100;
        Y = 4'b1010;
        // -------------------------------------
        // -------------  Current Time:  1900ns
        #100;
        Y = 4'b0110;
        // -------------------------------------
        // -------------  Current Time:  2000ns
        #100;
        Y = 4'b1111;
    end

endmodule

