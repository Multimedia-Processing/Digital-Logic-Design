module BUF_GATE (c, a);

input a;
output c;

    buf(c, a);

endmodule