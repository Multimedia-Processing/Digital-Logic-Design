module BUF_GATE_A (c, a);

input a;
output c;

    buf(c, a);

endmodule