
`timescale 1ns/1ps

module T;
    reg [7:0] D = 8'b01011111;
    wire Zero;
    wire One;


    all_zero_one UUT (
        .D(D),
        .Zero(Zero),
        .One(One));

    initial
    begin
      #1000 // Final time:  1000 ns
        $stop;
    end

    initial begin
        // -------------  Current Time:  100ns
        #100;
        D = 8'b11001000;
        // -------------------------------------
        // -------------  Current Time:  200ns
        #100;
        D = 8'b00000000;
        // -------------------------------------
        // -------------  Current Time:  300ns
        #100;
        D = 8'b00011101;
        // -------------------------------------
        // -------------  Current Time:  400ns
        #100;
        D = 8'b11101010;
        // -------------------------------------
        // -------------  Current Time:  500ns
        #100;
        D = 8'b01110011;
        // -------------------------------------
        // -------------  Current Time:  600ns
        #100;
        D = 8'b11111111;
        // -------------------------------------
        // -------------  Current Time:  700ns
        #100;
        D = 8'b10101000;
        // -------------------------------------
        // -------------  Current Time:  800ns
        #100;
        D = 8'b00111111;
        // -------------------------------------
        // -------------  Current Time:  900ns
        #100;
        D = 8'b01100110;
        // -------------------------------------
        // -------------  Current Time:  1000ns
        #100;
        CHECK_Zero(1'b0);
        D = 8'b11001000;
    end

endmodule

