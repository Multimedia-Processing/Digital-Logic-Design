module traffic_lights ();

endmodule // traffic_lights
