
`timescale 1ns/1ps

module T;
    reg I = 1'b0;
    reg C = 1'b1;
    wire O1;
    wire O2;
    wire O3;


    tri_gate UUT (
        .I(I),
        .C(C),
        .O1(O1),
        .O2(O2),
        .O3(O3));

    initial
    begin
      #1000 // Final time:  1000 ns
        $stop;
    end

    initial begin
        // -------------  Current Time:  100ns
        #100;
        I = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  200ns
        #100;
        I = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  300ns
        #100;
        I = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  400ns
        #100;
        I = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  500ns
        #100;
        I = 1'b1;
        C = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  600ns
        #100;
        I = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  700ns
        #100;
        I = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  800ns
        #100;
        I = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  900ns
        #100;
        I = 1'b1;
    end

endmodule

