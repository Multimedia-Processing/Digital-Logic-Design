module buf_gate (A,C);
    input A;
    output C;
    
    buf(C,A);
    
endmodule