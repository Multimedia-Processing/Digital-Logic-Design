module snake (clock, reset, turn, display);

endmodule // snake
