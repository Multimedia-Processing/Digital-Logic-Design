module up_counter_seven_segment_display ();

endmodule // up_counter_seven_segment_display
