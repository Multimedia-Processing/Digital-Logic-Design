module buf_gate (a, c);

  input a ;
  output c ;

  buf (c, a);

endmodule // buf_gate
