module nor_gate (a, b, c);

  input a, b ;
  output c ;

  nor (c, a, b);

endmodule // nor_gate
