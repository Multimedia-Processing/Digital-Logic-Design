// Ch02 and_gate.v
// �G��J�ιh (�h�h�y�z)

module and_gate (A, B, O);
input  A, B;	// A, B �@�줸��J
output O;	// O    �@�줸��X

and (O, A, B);

endmodule
